module mgmt_core ( VPWR, VGND, core_clk, flash_cs_n, flash_clk, flash_io0_oeb, 
        flash_io1_oeb, flash_io2_oeb, flash_io3_oeb, flash_io0_do, 
        flash_io1_do, flash_io2_do, flash_io3_do, flash_io0_di, flash_io1_di, 
        flash_io2_di, flash_io3_di, spi_clk, spi_cs_n, spi_mosi, spi_miso, 
        spi_sdoenb, mprj_wb_iena, mprj_cyc_o, mprj_stb_o, mprj_we_o, 
        mprj_sel_o, mprj_adr_o, mprj_dat_o, mprj_dat_i, mprj_ack_i, hk_dat_i, 
        hk_stb_o, hk_cyc_o, hk_ack_i, serial_tx, serial_rx, debug_in, 
        debug_out, debug_oeb, debug_mode, uart_enabled, gpio_out_pad, 
        gpio_in_pad, gpio_inenb_pad, gpio_mode0_pad, gpio_mode1_pad, la_output, 
        la_input, la_oenb, la_iena, qspi_enabled, spi_enabled, trap, 
        user_irq_ena, user_irq, clk_in, clk_out, resetn_in, resetn_out, 
        serial_load_in, serial_load_out, serial_data_2_in, serial_data_2_out, 
        serial_resetn_in, serial_resetn_out, serial_clock_in, serial_clock_out, 
        rstb_l_in, rstb_l_out, por_l_in, por_l_out, porb_h_in, porb_h_out, 
        gpio_outenb_pad_BAR, core_rstn_BAR );
  output [3:0] mprj_sel_o;
  output [31:0] mprj_adr_o;
  output [31:0] mprj_dat_o;
  input [31:0] mprj_dat_i;
  input [31:0] hk_dat_i;
  output [127:0] la_output;
  input [127:0] la_input;
  output [127:0] la_oenb;
  output [127:0] la_iena;
  output [2:0] user_irq_ena;
  input [5:0] user_irq;
  input core_clk, flash_io0_di, flash_io1_di, flash_io2_di, flash_io3_di,
         spi_miso, mprj_ack_i, hk_ack_i, serial_rx, debug_in, gpio_in_pad,
         clk_in, resetn_in, serial_load_in, serial_data_2_in, serial_resetn_in,
         serial_clock_in, rstb_l_in, por_l_in, porb_h_in, core_rstn_BAR;
  output flash_cs_n, flash_clk, flash_io0_oeb, flash_io1_oeb, flash_io2_oeb,
         flash_io3_oeb, flash_io0_do, flash_io1_do, flash_io2_do, flash_io3_do,
         spi_clk, spi_cs_n, spi_mosi, spi_sdoenb, mprj_wb_iena, mprj_cyc_o,
         mprj_stb_o, mprj_we_o, hk_stb_o, hk_cyc_o, serial_tx, debug_out,
         debug_oeb, debug_mode, uart_enabled, gpio_out_pad, gpio_inenb_pad,
         gpio_mode0_pad, gpio_mode1_pad, qspi_enabled, spi_enabled, trap,
         clk_out, resetn_out, serial_load_out, serial_data_2_out,
         serial_resetn_out, serial_clock_out, rstb_l_out, por_l_out,
         porb_h_out, gpio_outenb_pad_BAR;
  inout VPWR,  VGND;
  wire   core_rstn, hk_stb_o, n6130, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n6131, n6132, n6133, sys_uart_rx, dbg_uart_dbg_uart_rx,
         dbg_uart_dbg_uart_tx, sys_uart_tx, uart_enabled_o, sys_rst,
         mgmtsoc_zero1, mgmtsoc_pending_re, mgmtsoc_pending_r, dff2_en,
         mgmtsoc_litespisdrphycore_dq_o, mgmtsoc_litespisdrphycore_clk,
         mgmtsoc_litespisdrphycore_posedge_reg2,
         mgmtsoc_port_master_user_port_sink_valid,
         \mgmtsoc_port_master_user_port_sink_payload_mask[0] ,
         \litespi_request[1] , litespi_tx_mux_sel,
         mgmtsoc_litespimmap_burst_cs, spi_master_loopback,
         rs232phy_rs232phytx_state, uart_phy_tx_tick, uart_phy_tx_sink_valid,
         rs232phy_rs232phyrx_state, uart_phy_rx_tick, uart_phy_rx_rx,
         uart_phy_rx_rx_d, uart_pending_re,
         uartwishbonebridge_rs232phytx_state, dbg_uart_tx_tick,
         uartwishbonebridge_rs232phyrx_state, dbg_uart_rx_tick, dbg_uart_rx_rx,
         dbg_uart_rx_rx_d, dbg_uart_incr, gpioin0_i01, gpioin0_pending_re,
         gpioin0_pending_r, gpioin1_i01, gpioin1_pending_re, gpioin1_pending_r,
         gpioin2_i01, gpioin2_pending_re, gpioin2_pending_r,
         gpioin3_gpioin3_in_pads_n_d, gpioin3_i01, gpioin3_pending_re,
         gpioin3_pending_r, gpioin4_gpioin4_in_pads_n_d, gpioin4_i01,
         gpioin4_pending_re, gpioin4_pending_r, gpioin5_gpioin5_in_pads_n_d,
         gpioin5_i01, gpioin5_pending_re, gpioin5_pending_r, state,
         mgmtsoc_ibus_ibus_ack, mgmtsoc_dbus_dbus_ack,
         mgmtsoc_vexriscv_debug_bus_ack, dff_bus_ack, dff2_bus_ack,
         mgmtsoc_reset_re, \mgmtsoc_master_status_status[1] , csrbank5_ien0_w,
         csrbank5_oe0_w, csrbank5_in_w, spi_master_control_re, csrbank10_en0_w,
         csrbank10_update_value0_w, mgmtsoc_zero2, \uart_status_status[1] ,
         csrbank13_mode0_w, csrbank13_edge0_w, gpioin0_i02, csrbank14_mode0_w,
         csrbank14_edge0_w, gpioin1_i02, csrbank15_mode0_w, csrbank15_edge0_w,
         gpioin2_i02, csrbank16_in_w, csrbank16_mode0_w, csrbank16_edge0_w,
         gpioin3_i02, csrbank17_in_w, csrbank17_mode0_w, csrbank17_edge0_w,
         gpioin4_i02, csrbank18_in_w, csrbank18_mode0_w, csrbank18_edge0_w,
         gpioin5_i02, \interface1_bank_bus_dat_r[0] ,
         \interface2_bank_bus_dat_r[0] , \interface5_bank_bus_dat_r[0] ,
         \interface7_bank_bus_dat_r[0] , \interface8_bank_bus_dat_r[0] ,
         \interface12_bank_bus_dat_r[0] , \interface13_bank_bus_dat_r[0] ,
         \interface14_bank_bus_dat_r[0] , \interface15_bank_bus_dat_r[0] ,
         \interface16_bank_bus_dat_r[0] , \interface17_bank_bus_dat_r[0] ,
         \interface18_bank_bus_dat_r[0] , mgmtsoc_dbus_dbus_we,
         \mgmtsoc_litespisdrphycore_dq_i[1] ,
         mgmtsoc_vexriscv_transfer_complete,
         mgmtsoc_vexriscv_transfer_wait_for_ack, mgmtsoc_vexriscv_o_cmd_ready,
         mgmtsoc_vexriscv_o_resetOut, mgmtsoc_update_value_re,
         mgmtsoc_vexriscv_reset_debug_logic, mgmtsoc_vexriscv_debug_reset,
         mgmtsoc_vexriscv_i_cmd_payload_wr, mgmtsoc_vexriscv_i_cmd_valid,
         mgmtsoc_zero_trigger_d, mgmtsoc_litespisdrphycore_posedge_reg, N3577,
         N3578, N3579, N3580, N3581, N3582, N3583, N3584, N3585, N3586, N3587,
         N3588, N3589, N3590, N3591, N3592, N3593, N3594, N3595, N3596, N3597,
         N3598, N3599, N3600, N3601, N3602, N3603, N3644, N3645, N3646, N3647,
         N3648, N3649, N3650, N3651, N3652, N3653, N3654, N3655, N3656, N3657,
         N3658, N3659, N3660, N3661, N3662, N3663, N3664, N3665, N3666, N3667,
         N3668, N3669, N3670, uart_tx_trigger_d, uart_rx_trigger_d,
         gpioin0_gpioin0_trigger_d, gpioin1_gpioin1_trigger_d,
         gpioin2_gpioin2_trigger_d, gpioin3_gpioin3_trigger_d,
         gpioin4_gpioin4_trigger_d, gpioin5_gpioin5_trigger_d, N4099, N4100,
         N4101, N4102, N4103, N4104, N4105, N4106, N4107, N4108, N4109, N4110,
         N4111, N4112, N4113, N4114, N4115, N4116, N4117, N4118, N4119, N4120,
         N4121, N4122, N4123, N4124, N4125, N4126, N4127, N4128, N4129, N4130,
         N4141, N4152, N4243, N4244, N4245, N4246, N4247, N4248, N4249, N4250,
         N4251, N4252, N4253, N4254, N4255, N4256, N4257, N4258, N4259, N4260,
         N4261, N4262, N4263, N4264, N4265, N4266, N4267, N4268, N4269, N4270,
         N4271, N4272, N4273, N4274, N4292, N4293, N4294, N4295, N4296, N4297,
         N4298, N4299, N4331, N4463, N4464, N4465, N4466, N4467, N4468, N4469,
         N4470, N4471, N4472, N4473, N4474, N4475, N4476, N4477, N4478, N4479,
         N4480, N4481, N4482, N4483, N4484, N4485, N4486, N4487, N4488, N4489,
         N4490, N4491, N4492, N4493, N4494, N4505, N4516, N4585, N4586, N4587,
         N4588, N4589, N4590, N4591, N4592, N4593, N4594, N4595, N4596, N4597,
         N4598, N4599, N4600, N4601, N4694, N4695, N4696, N4697, N4698, N4699,
         N4700, N4701, N4702, N4703, N4704, N4705, N4706, N4707, N4708, N4709,
         N4710, N4711, N4712, N4713, N4714, N4715, N4716, N4717, N4718, N4719,
         N4720, N4721, N4722, N4723, N4724, N4725, N4772, N4773, N4774, N4775,
         N4776, N4777, N4778, N4779, N4790, N4822, N4854, N4886, N4918, N4950,
         N4982, N4995, N4996, N4997, N5014, N5015, N5016, N5017, N5018, N5019,
         N5020, N5021, N5022, N5023, N5024, N5025, N5026, N5027, N5028, N5029,
         N5030, N5031, N5032, N5033, N5034, N5035, N5036, N5037, N5038, N5039,
         N5040, N5041, N5042, N5043, N5044, N5045, N5046, N5047, N5048, N5049,
         N5050, N5051, N5052, N5053, N5054, N5055, N5056, N5057, N5058, N5059,
         N5060, N5061, N5062, N5063, N5064, N5065, N5066, N5067, N5068, N5069,
         N5070, N5071, N5072, N5073, N5074, N5075, N5076, N5077, N5168, N5235,
         N5281, N5358, N5394, N5395, N5400, N5401, N5402, N5403, N5404, N5405,
         N5406, N5407, N5408, N5409, N5410, N5411, N5412, N5413, N5414, N5415,
         N5416, N5417, N5418, N5419, N5420, N5421, N5422, N5423, N5424, N5425,
         N5426, N5427, N5428, N5429, N5430, N5431, N5432, N5433, N5443, N5444,
         N5445, N5446, N5447, N5448, N5449, N5450, N5453, N5454, N5589, N5618,
         N5643, N5644, N5645, N5646, N5647, N5648, N5649, N5650, N5651, N5652,
         N5653, N5654, N5655, N5656, N5657, N5658, N5702, N5703, N5704, N5707,
         N5710, N5711, N5756, N5757, N5758, N6207, N6215, N6223, N6228, N6231,
         N6236, N6239, N6244, N6247, N6248, N6249, N6252, N6253, N6254, N6255,
         N6262, N6263, N6264, N6265, N6270, N6275, N6280, N6285, N6290, N6298,
         N6299, N6300, N6301, N6302, N6303, N6304, N6326, multiregimpl0_regs0,
         multiregimpl1_regs0, multiregimpl2_regs0, multiregimpl134_regs0,
         multiregimpl135_regs0, multiregimpl136_regs0, \storage[0][7] ,
         \storage[0][6] , \storage[0][5] , \storage[0][4] , \storage[0][3] ,
         \storage[0][2] , \storage[0][1] , \storage[0][0] , \storage[1][7] ,
         \storage[1][6] , \storage[1][5] , \storage[1][4] , \storage[1][3] ,
         \storage[1][2] , \storage[1][1] , \storage[1][0] , \storage[2][7] ,
         \storage[2][6] , \storage[2][5] , \storage[2][4] , \storage[2][3] ,
         \storage[2][2] , \storage[2][1] , \storage[2][0] , \storage[3][7] ,
         \storage[3][6] , \storage[3][5] , \storage[3][4] , \storage[3][3] ,
         \storage[3][2] , \storage[3][1] , \storage[3][0] , \storage[4][7] ,
         \storage[4][6] , \storage[4][5] , \storage[4][4] , \storage[4][3] ,
         \storage[4][2] , \storage[4][1] , \storage[4][0] , \storage[5][7] ,
         \storage[5][6] , \storage[5][5] , \storage[5][4] , \storage[5][3] ,
         \storage[5][2] , \storage[5][1] , \storage[5][0] , \storage[6][7] ,
         \storage[6][6] , \storage[6][5] , \storage[6][4] , \storage[6][3] ,
         \storage[6][2] , \storage[6][1] , \storage[6][0] , \storage[7][7] ,
         \storage[7][6] , \storage[7][5] , \storage[7][4] , \storage[7][3] ,
         \storage[7][2] , \storage[7][1] , \storage[7][0] , \storage[8][7] ,
         \storage[8][6] , \storage[8][5] , \storage[8][4] , \storage[8][3] ,
         \storage[8][2] , \storage[8][1] , \storage[8][0] , \storage[9][7] ,
         \storage[9][6] , \storage[9][5] , \storage[9][4] , \storage[9][3] ,
         \storage[9][2] , \storage[9][1] , \storage[9][0] , \storage[10][7] ,
         \storage[10][6] , \storage[10][5] , \storage[10][4] ,
         \storage[10][3] , \storage[10][2] , \storage[10][1] ,
         \storage[10][0] , \storage[11][7] , \storage[11][6] ,
         \storage[11][5] , \storage[11][4] , \storage[11][3] ,
         \storage[11][2] , \storage[11][1] , \storage[11][0] ,
         \storage[12][7] , \storage[12][6] , \storage[12][5] ,
         \storage[12][4] , \storage[12][3] , \storage[12][2] ,
         \storage[12][1] , \storage[12][0] , \storage[13][7] ,
         \storage[13][6] , \storage[13][5] , \storage[13][4] ,
         \storage[13][3] , \storage[13][2] , \storage[13][1] ,
         \storage[13][0] , \storage[14][7] , \storage[14][6] ,
         \storage[14][5] , \storage[14][4] , \storage[14][3] ,
         \storage[14][2] , \storage[14][1] , \storage[14][0] ,
         \storage[15][7] , \storage[15][6] , \storage[15][5] ,
         \storage[15][4] , \storage[15][3] , \storage[15][2] ,
         \storage[15][1] , \storage[15][0] , \storage_1[0][7] ,
         \storage_1[0][6] , \storage_1[0][5] , \storage_1[0][4] ,
         \storage_1[0][3] , \storage_1[0][2] , \storage_1[0][1] ,
         \storage_1[0][0] , \storage_1[1][7] , \storage_1[1][6] ,
         \storage_1[1][5] , \storage_1[1][4] , \storage_1[1][3] ,
         \storage_1[1][2] , \storage_1[1][1] , \storage_1[1][0] ,
         \storage_1[2][7] , \storage_1[2][6] , \storage_1[2][5] ,
         \storage_1[2][4] , \storage_1[2][3] , \storage_1[2][2] ,
         \storage_1[2][1] , \storage_1[2][0] , \storage_1[3][7] ,
         \storage_1[3][6] , \storage_1[3][5] , \storage_1[3][4] ,
         \storage_1[3][3] , \storage_1[3][2] , \storage_1[3][1] ,
         \storage_1[3][0] , \storage_1[4][7] , \storage_1[4][6] ,
         \storage_1[4][5] , \storage_1[4][4] , \storage_1[4][3] ,
         \storage_1[4][2] , \storage_1[4][1] , \storage_1[4][0] ,
         \storage_1[5][7] , \storage_1[5][6] , \storage_1[5][5] ,
         \storage_1[5][4] , \storage_1[5][3] , \storage_1[5][2] ,
         \storage_1[5][1] , \storage_1[5][0] , \storage_1[6][7] ,
         \storage_1[6][6] , \storage_1[6][5] , \storage_1[6][4] ,
         \storage_1[6][3] , \storage_1[6][2] , \storage_1[6][1] ,
         \storage_1[6][0] , \storage_1[7][7] , \storage_1[7][6] ,
         \storage_1[7][5] , \storage_1[7][4] , \storage_1[7][3] ,
         \storage_1[7][2] , \storage_1[7][1] , \storage_1[7][0] ,
         \storage_1[8][7] , \storage_1[8][6] , \storage_1[8][5] ,
         \storage_1[8][4] , \storage_1[8][3] , \storage_1[8][2] ,
         \storage_1[8][1] , \storage_1[8][0] , \storage_1[9][7] ,
         \storage_1[9][6] , \storage_1[9][5] , \storage_1[9][4] ,
         \storage_1[9][3] , \storage_1[9][2] , \storage_1[9][1] ,
         \storage_1[9][0] , \storage_1[10][7] , \storage_1[10][6] ,
         \storage_1[10][5] , \storage_1[10][4] , \storage_1[10][3] ,
         \storage_1[10][2] , \storage_1[10][1] , \storage_1[10][0] ,
         \storage_1[11][7] , \storage_1[11][6] , \storage_1[11][5] ,
         \storage_1[11][4] , \storage_1[11][3] , \storage_1[11][2] ,
         \storage_1[11][1] , \storage_1[11][0] , \storage_1[12][7] ,
         \storage_1[12][6] , \storage_1[12][5] , \storage_1[12][4] ,
         \storage_1[12][3] , \storage_1[12][2] , \storage_1[12][1] ,
         \storage_1[12][0] , \storage_1[13][7] , \storage_1[13][6] ,
         \storage_1[13][5] , \storage_1[13][4] , \storage_1[13][3] ,
         \storage_1[13][2] , \storage_1[13][1] , \storage_1[13][0] ,
         \storage_1[14][7] , \storage_1[14][6] , \storage_1[14][5] ,
         \storage_1[14][4] , \storage_1[14][3] , \storage_1[14][2] ,
         \storage_1[14][1] , \storage_1[14][0] , \storage_1[15][7] ,
         \storage_1[15][6] , \storage_1[15][5] , \storage_1[15][4] ,
         \storage_1[15][3] , \storage_1[15][2] , \storage_1[15][1] ,
         \storage_1[15][0] , _2_net_, \RAM256/Do0_pre[1][31] ,
         \RAM256/Do0_pre[1][30] , \RAM256/Do0_pre[1][29] ,
         \RAM256/Do0_pre[1][28] , \RAM256/Do0_pre[1][27] ,
         \RAM256/Do0_pre[1][26] , \RAM256/Do0_pre[1][25] ,
         \RAM256/Do0_pre[1][24] , \RAM256/Do0_pre[1][23] ,
         \RAM256/Do0_pre[1][22] , \RAM256/Do0_pre[1][21] ,
         \RAM256/Do0_pre[1][20] , \RAM256/Do0_pre[1][19] ,
         \RAM256/Do0_pre[1][18] , \RAM256/Do0_pre[1][17] ,
         \RAM256/Do0_pre[1][16] , \RAM256/Do0_pre[1][15] ,
         \RAM256/Do0_pre[1][14] , \RAM256/Do0_pre[1][13] ,
         \RAM256/Do0_pre[1][12] , \RAM256/Do0_pre[1][11] ,
         \RAM256/Do0_pre[1][10] , \RAM256/Do0_pre[1][9] ,
         \RAM256/Do0_pre[1][8] , \RAM256/Do0_pre[1][7] ,
         \RAM256/Do0_pre[1][6] , \RAM256/Do0_pre[1][5] ,
         \RAM256/Do0_pre[1][4] , \RAM256/Do0_pre[1][3] ,
         \RAM256/Do0_pre[1][2] , \RAM256/Do0_pre[1][1] ,
         \RAM256/Do0_pre[1][0] , \RAM256/Do0_pre[0][31] ,
         \RAM256/Do0_pre[0][30] , \RAM256/Do0_pre[0][29] ,
         \RAM256/Do0_pre[0][28] , \RAM256/Do0_pre[0][27] ,
         \RAM256/Do0_pre[0][26] , \RAM256/Do0_pre[0][25] ,
         \RAM256/Do0_pre[0][24] , \RAM256/Do0_pre[0][23] ,
         \RAM256/Do0_pre[0][22] , \RAM256/Do0_pre[0][21] ,
         \RAM256/Do0_pre[0][20] , \RAM256/Do0_pre[0][19] ,
         \RAM256/Do0_pre[0][18] , \RAM256/Do0_pre[0][17] ,
         \RAM256/Do0_pre[0][16] , \RAM256/Do0_pre[0][15] ,
         \RAM256/Do0_pre[0][14] , \RAM256/Do0_pre[0][13] ,
         \RAM256/Do0_pre[0][12] , \RAM256/Do0_pre[0][11] ,
         \RAM256/Do0_pre[0][10] , \RAM256/Do0_pre[0][9] ,
         \RAM256/Do0_pre[0][8] , \RAM256/Do0_pre[0][7] ,
         \RAM256/Do0_pre[0][6] , \RAM256/Do0_pre[0][5] ,
         \RAM256/Do0_pre[0][4] , \RAM256/Do0_pre[0][3] ,
         \RAM256/Do0_pre[0][2] , \RAM256/Do0_pre[0][1] ,
         \RAM256/Do0_pre[0][0] , \RAM256/SEL0[1] , \RAM256/SEL0[0] ,
         \RAM256/VGND , \RAM256/VPWR , n3088, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n266, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3089, n3118, n3119, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129;
  wire   [7:0] mgmtsoc_interrupt;
  wire   [31:0] mgmtsoc_bus_errors_status;
  wire   [31:0] mgmtsoc_value;
  wire   [3:0] dff_we;
  wire   [3:0] dff2_we;
  wire   [31:0] dff2_bus_dat_r;
  wire   [7:0] mgmtsoc_litespisdrphycore_div;
  wire   [31:0] mgmtsoc_litespisdrphycore_sr_out;
  wire   [31:0] mgmtsoc_litespisdrphycore_source_payload_data;
  wire   [7:0] mgmtsoc_litespisdrphycore_cnt;
  wire   [3:0] mgmtsoc_litespisdrphycore_count;
  wire   [1:0] litespiphy_state;
  wire   [7:0] mgmtsoc_litespisdrphycore_sr_cnt;
  wire   [31:0] mgmtsoc_port_master_user_port_sink_payload_data;
  wire   [5:0] mgmtsoc_port_master_user_port_sink_payload_len;
  wire   [3:0] mgmtsoc_port_master_user_port_sink_payload_width;
  wire   [7:0] mgmtsoc_litespimmap_spi_dummy_bits;
  wire   [8:0] mgmtsoc_litespimmap_count;
  wire   [3:0] litespi_state;
  wire   [29:0] mgmtsoc_litespimmap_burst_adr;
  wire   [7:6] mgmtsoc_master_len;
  wire   [5:0] mgmtsoc_master_tx_fifo_sink_payload_len;
  wire   [3:0] mgmtsoc_master_tx_fifo_sink_payload_width;
  wire   [7:0] mgmtsoc_master_tx_fifo_sink_payload_mask;
  wire   [31:0] mgmtsoc_master_rxtx_w;
  wire   [7:0] spi_master_length0;
  wire   [7:0] spi_master_mosi;
  wire   [7:0] spi_master_miso_status;
  wire   [15:0] spi_master_clk_divider1;
  wire   [15:0] spi_master_clk_divider0;
  wire   [1:0] spimaster_state;
  wire   [2:0] spi_master_count;
  wire   [3:0] uart_phy_tx_count;
  wire   [7:0] uart_phy_tx_data;
  wire   [3:0] uart_phy_rx_count;
  wire   [7:0] uart_phy_rx_data;
  wire   [1:0] uart_pending_r;
  wire   [1:0] uart_pending_status;
  wire   [7:0] uart_tx_fifo_fifo_out_payload_data;
  wire   [4:0] uart_tx_fifo_level0;
  wire   [3:0] uart_tx_fifo_produce;
  wire   [3:0] uart_tx_fifo_rdport_adr;
  wire   [7:0] uart_rx_fifo_fifo_out_payload_data;
  wire   [4:0] uart_rx_fifo_level0;
  wire   [3:0] uart_rx_fifo_produce;
  wire   [3:0] uart_rx_fifo_rdport_adr;
  wire   [29:0] dbg_uart_wishbone_adr;
  wire   [31:0] dbg_uart_wishbone_dat_w;
  wire   [1:0] dbg_uart_bytes_count;
  wire   [7:0] dbg_uart_words_count;
  wire   [7:0] dbg_uart_length;
  wire   [3:0] dbg_uart_tx_count;
  wire   [7:0] dbg_uart_tx_data;
  wire   [3:0] dbg_uart_rx_count;
  wire   [7:0] dbg_uart_rx_data;
  wire   [2:0] uartwishbonebridge_state;
  wire   [7:0] dbg_uart_cmd;
  wire   [19:0] dbg_uart_count;
  wire   [31:0] mgmtsoc_ibus_ibus_dat_r;
  wire   [1:0] grant;
  wire   [2:0] request;
  wire   [6:0] slave_sel_r;
  wire   [31:0] mgmtsoc_vexriscv_debug_bus_dat_r;
  wire   [19:0] count;
  wire   [1:0] csrbank0_reset0_w;
  wire   [31:0] csrbank0_scratch0_w;
  wire   [15:12] csrbank3_master_phyconfig0_w;
  wire   [31:0] csrbank6_ien3_w;
  wire   [31:0] csrbank6_ien2_w;
  wire   [31:0] csrbank6_ien1_w;
  wire   [31:0] csrbank6_ien0_w;
  wire   [31:0] csrbank6_oe3_w;
  wire   [31:0] csrbank6_oe2_w;
  wire   [31:0] csrbank6_oe1_w;
  wire   [31:0] csrbank6_oe0_w;
  wire   [7:0] csrbank9_control0_w;
  wire   [16:0] csrbank9_cs0_w;
  wire   [31:0] csrbank10_load0_w;
  wire   [31:0] csrbank10_reload0_w;
  wire   [31:0] csrbank10_value_w;
  wire   [1:0] csrbank11_ev_enable0_w;
  wire   [31:0] interface0_bank_bus_dat_r;
  wire   [31:0] interface3_bank_bus_dat_r;
  wire   [31:0] interface4_bank_bus_dat_r;
  wire   [31:0] interface6_bank_bus_dat_r;
  wire   [31:0] interface9_bank_bus_dat_r;
  wire   [31:0] interface10_bank_bus_dat_r;
  wire   [31:0] interface11_bank_bus_dat_r;
  wire   [31:0] interface19_bank_bus_dat_r;
  wire   [29:0] mgmtsoc_ibus_ibus_adr;
  wire   [29:0] mgmtsoc_dbus_dbus_adr;
  wire   [31:0] mgmtsoc_dbus_dbus_dat_w;
  wire   [3:0] mgmtsoc_dbus_dbus_sel;
  wire   [7:0] spi_master_mosi_data;
  wire   [2:0] spi_master_mosi_sel;
  wire   [7:0] spi_master_miso_data;
  wire   [31:0] mgmtsoc_vexriscv_o_rsp_data;
  wire   [31:0] mgmtsoc_vexriscv_i_cmd_payload_data;
  wire   [7:0] mgmtsoc_vexriscv_i_cmd_payload_address;
  wire   [31:0] uart_phy_tx_phase;
  wire   [31:0] uart_phy_rx_phase;
  wire   [31:0] dbg_uart_tx_phase;
  wire   [31:0] dbg_uart_rx_phase;
  assign core_rstn = core_rstn_BAR;
  assign mprj_stb_o = hk_stb_o;
  assign gpio_outenb_pad_BAR = csrbank5_oe0_w;

  RAM128 RAM128 ( .CLK(n6106), .EN0(dff2_en), .VGND(1'b0), .VPWR(1'b0), .A0(
        mprj_adr_o[8:2]), .Di0(mprj_dat_o), .Do0(dff2_bus_dat_r), .WE0(dff2_we) );
  VexRiscv VexRiscv ( .vccd1(VPWR), .vssd1(VGND), .externalResetVector({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .timerInterrupt(1'b0), 
        .softwareInterrupt(1'b0), .externalInterruptArray({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        mgmtsoc_interrupt}), .debug_bus_cmd_valid(mgmtsoc_vexriscv_i_cmd_valid), .debug_bus_cmd_ready(mgmtsoc_vexriscv_o_cmd_ready), 
        .debug_bus_cmd_payload_wr(mgmtsoc_vexriscv_i_cmd_payload_wr), 
        .debug_bus_cmd_payload_address({
        mgmtsoc_vexriscv_i_cmd_payload_address[7:2], 1'b0, 1'b0}), 
        .debug_bus_cmd_payload_data(mgmtsoc_vexriscv_i_cmd_payload_data), 
        .debug_bus_rsp_data(mgmtsoc_vexriscv_o_rsp_data), .debug_resetOut(
        mgmtsoc_vexriscv_o_resetOut), .iBusWishbone_CYC(request[0]), 
        .iBusWishbone_ACK(mgmtsoc_ibus_ibus_ack), .iBusWishbone_DAT_MISO(
        mgmtsoc_ibus_ibus_dat_r), .iBusWishbone_ERR(1'b0), .dBusWishbone_CYC(
        request[1]), .dBusWishbone_ACK(mgmtsoc_dbus_dbus_ack), 
        .dBusWishbone_WE(mgmtsoc_dbus_dbus_we), .dBusWishbone_ADR(
        mgmtsoc_dbus_dbus_adr), .dBusWishbone_DAT_MISO({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .dBusWishbone_DAT_MOSI(
        mgmtsoc_dbus_dbus_dat_w), .dBusWishbone_SEL(mgmtsoc_dbus_dbus_sel), 
        .dBusWishbone_ERR(1'b0), .clk(n6111), .reset(_2_net_), .debugReset(
        sys_rst), .\iBusWishbone_ADR[29] (mgmtsoc_ibus_ibus_adr[29]), 
        .\iBusWishbone_ADR[28] (mgmtsoc_ibus_ibus_adr[28]), 
        .\iBusWishbone_ADR[27] (mgmtsoc_ibus_ibus_adr[27]), 
        .\iBusWishbone_ADR[26] (mgmtsoc_ibus_ibus_adr[26]), 
        .\iBusWishbone_ADR[25] (mgmtsoc_ibus_ibus_adr[25]), 
        .\iBusWishbone_ADR[24] (mgmtsoc_ibus_ibus_adr[24]), 
        .\iBusWishbone_ADR[23] (mgmtsoc_ibus_ibus_adr[23]), 
        .\iBusWishbone_ADR[22] (mgmtsoc_ibus_ibus_adr[22]), 
        .\iBusWishbone_ADR[21] (mgmtsoc_ibus_ibus_adr[21]), 
        .\iBusWishbone_ADR[20] (mgmtsoc_ibus_ibus_adr[20]), 
        .\iBusWishbone_ADR[19] (mgmtsoc_ibus_ibus_adr[19]), 
        .\iBusWishbone_ADR[18] (mgmtsoc_ibus_ibus_adr[18]), 
        .\iBusWishbone_ADR[17] (mgmtsoc_ibus_ibus_adr[17]), 
        .\iBusWishbone_ADR[16] (mgmtsoc_ibus_ibus_adr[16]), 
        .\iBusWishbone_ADR[15] (mgmtsoc_ibus_ibus_adr[15]), 
        .\iBusWishbone_ADR[14] (mgmtsoc_ibus_ibus_adr[14]), 
        .\iBusWishbone_ADR[13] (mgmtsoc_ibus_ibus_adr[13]), 
        .\iBusWishbone_ADR[12] (mgmtsoc_ibus_ibus_adr[12]), 
        .\iBusWishbone_ADR[11] (mgmtsoc_ibus_ibus_adr[11]), 
        .\iBusWishbone_ADR[10] (mgmtsoc_ibus_ibus_adr[10]), 
        .\iBusWishbone_ADR[9] (mgmtsoc_ibus_ibus_adr[9]), 
        .\iBusWishbone_ADR[8] (mgmtsoc_ibus_ibus_adr[8]), 
        .\iBusWishbone_ADR[7] (mgmtsoc_ibus_ibus_adr[7]), 
        .\iBusWishbone_ADR[6] (mgmtsoc_ibus_ibus_adr[6]), 
        .\iBusWishbone_ADR[5] (mgmtsoc_ibus_ibus_adr[5]), 
        .\iBusWishbone_ADR[4] (mgmtsoc_ibus_ibus_adr[4]), 
        .\iBusWishbone_ADR[3]_BAR (mgmtsoc_ibus_ibus_adr[3]), 
        .\iBusWishbone_ADR[2] (mgmtsoc_ibus_ibus_adr[2]), 
        .\iBusWishbone_ADR[1] (mgmtsoc_ibus_ibus_adr[1]), 
        .\iBusWishbone_ADR[0] (mgmtsoc_ibus_ibus_adr[0]) );
  RAM128 \RAM256/BANK128[1].RAM128  ( .CLK(n6039), .EN0(\RAM256/SEL0[1] ), 
        .VGND(\RAM256/VGND ), .VPWR(\RAM256/VPWR ), .A0(mprj_adr_o[8:2]), 
        .Di0(mprj_dat_o), .Do0({\RAM256/Do0_pre[1][31] , 
        \RAM256/Do0_pre[1][30] , \RAM256/Do0_pre[1][29] , 
        \RAM256/Do0_pre[1][28] , \RAM256/Do0_pre[1][27] , 
        \RAM256/Do0_pre[1][26] , \RAM256/Do0_pre[1][25] , 
        \RAM256/Do0_pre[1][24] , \RAM256/Do0_pre[1][23] , 
        \RAM256/Do0_pre[1][22] , \RAM256/Do0_pre[1][21] , 
        \RAM256/Do0_pre[1][20] , \RAM256/Do0_pre[1][19] , 
        \RAM256/Do0_pre[1][18] , \RAM256/Do0_pre[1][17] , 
        \RAM256/Do0_pre[1][16] , \RAM256/Do0_pre[1][15] , 
        \RAM256/Do0_pre[1][14] , \RAM256/Do0_pre[1][13] , 
        \RAM256/Do0_pre[1][12] , \RAM256/Do0_pre[1][11] , 
        \RAM256/Do0_pre[1][10] , \RAM256/Do0_pre[1][9] , 
        \RAM256/Do0_pre[1][8] , \RAM256/Do0_pre[1][7] , \RAM256/Do0_pre[1][6] , 
        \RAM256/Do0_pre[1][5] , \RAM256/Do0_pre[1][4] , \RAM256/Do0_pre[1][3] , 
        \RAM256/Do0_pre[1][2] , \RAM256/Do0_pre[1][1] , \RAM256/Do0_pre[1][0] }), .WE0(dff_we) );
  RAM128 \RAM256/BANK128[0].RAM128  ( .CLK(n6105), .EN0(\RAM256/SEL0[0] ), 
        .VGND(\RAM256/VGND ), .VPWR(\RAM256/VPWR ), .A0(mprj_adr_o[8:2]), 
        .Di0(mprj_dat_o), .Do0({\RAM256/Do0_pre[0][31] , 
        \RAM256/Do0_pre[0][30] , \RAM256/Do0_pre[0][29] , 
        \RAM256/Do0_pre[0][28] , \RAM256/Do0_pre[0][27] , 
        \RAM256/Do0_pre[0][26] , \RAM256/Do0_pre[0][25] , 
        \RAM256/Do0_pre[0][24] , \RAM256/Do0_pre[0][23] , 
        \RAM256/Do0_pre[0][22] , \RAM256/Do0_pre[0][21] , 
        \RAM256/Do0_pre[0][20] , \RAM256/Do0_pre[0][19] , 
        \RAM256/Do0_pre[0][18] , \RAM256/Do0_pre[0][17] , 
        \RAM256/Do0_pre[0][16] , \RAM256/Do0_pre[0][15] , 
        \RAM256/Do0_pre[0][14] , \RAM256/Do0_pre[0][13] , 
        \RAM256/Do0_pre[0][12] , \RAM256/Do0_pre[0][11] , 
        \RAM256/Do0_pre[0][10] , \RAM256/Do0_pre[0][9] , 
        \RAM256/Do0_pre[0][8] , \RAM256/Do0_pre[0][7] , \RAM256/Do0_pre[0][6] , 
        \RAM256/Do0_pre[0][5] , \RAM256/Do0_pre[0][4] , \RAM256/Do0_pre[0][3] , 
        \RAM256/Do0_pre[0][2] , \RAM256/Do0_pre[0][1] , \RAM256/Do0_pre[0][0] }), .WE0(dff_we) );
  dfnrq1 int_rst_reg ( .D(core_rstn), .CP(n6067), .Q(sys_rst) );
  dfnrq1 \mgmtsoc_litespisdrphycore_dq_i_reg[1]  ( .D(flash_io1_di), .CP(n6128), .Q(\mgmtsoc_litespisdrphycore_dq_i[1] ) );
  dfnrq1 multiregimpl134_regs0_reg ( .D(user_irq[3]), .CP(n6060), .Q(
        multiregimpl134_regs0) );
  dfnrq1 multiregimpl135_regs0_reg ( .D(user_irq[4]), .CP(n6053), .Q(
        multiregimpl135_regs0) );
  dfnrq1 multiregimpl136_regs0_reg ( .D(user_irq[5]), .CP(n6050), .Q(
        multiregimpl136_regs0) );
  dfnrq1 multiregimpl136_regs1_reg ( .D(multiregimpl136_regs0), .CP(n6050), 
        .Q(csrbank18_in_w) );
  dfnrq1 multiregimpl135_regs1_reg ( .D(multiregimpl135_regs0), .CP(n6050), 
        .Q(csrbank17_in_w) );
  dfnrq1 multiregimpl134_regs1_reg ( .D(multiregimpl134_regs0), .CP(n6050), 
        .Q(csrbank16_in_w) );
  dfnrq1 \spi_master_clk_divider1_reg[15]  ( .D(N5658), .CP(n6051), .Q(
        spi_master_clk_divider1[15]) );
  dfnrq1 \spi_master_clk_divider1_reg[14]  ( .D(N5657), .CP(n6051), .Q(
        spi_master_clk_divider1[14]) );
  dfnrq1 \spi_master_clk_divider1_reg[13]  ( .D(N5656), .CP(n6051), .Q(
        spi_master_clk_divider1[13]) );
  dfnrq1 \spi_master_clk_divider1_reg[12]  ( .D(N5655), .CP(n6051), .Q(
        spi_master_clk_divider1[12]) );
  dfnrq1 \spi_master_clk_divider1_reg[11]  ( .D(N5654), .CP(n6051), .Q(
        spi_master_clk_divider1[11]) );
  dfnrq1 \spi_master_clk_divider1_reg[10]  ( .D(N5653), .CP(n6051), .Q(
        spi_master_clk_divider1[10]) );
  dfnrq1 \spi_master_clk_divider1_reg[9]  ( .D(N5652), .CP(n6051), .Q(
        spi_master_clk_divider1[9]) );
  dfnrq1 \spi_master_clk_divider1_reg[8]  ( .D(N5651), .CP(n6051), .Q(
        spi_master_clk_divider1[8]) );
  dfnrq1 \spi_master_clk_divider1_reg[7]  ( .D(N5650), .CP(n6113), .Q(
        spi_master_clk_divider1[7]) );
  dfnrq1 \spi_master_clk_divider1_reg[6]  ( .D(N5649), .CP(n6027), .Q(
        spi_master_clk_divider1[6]) );
  dfnrq1 \spi_master_clk_divider1_reg[5]  ( .D(N5648), .CP(n6049), .Q(
        spi_master_clk_divider1[5]) );
  dfnrq1 \spi_master_clk_divider1_reg[4]  ( .D(N5647), .CP(n6027), .Q(
        spi_master_clk_divider1[4]) );
  dfnrq1 \spi_master_clk_divider1_reg[3]  ( .D(N5646), .CP(n6043), .Q(
        spi_master_clk_divider1[3]) );
  dfnrq1 \spi_master_clk_divider1_reg[2]  ( .D(N5645), .CP(n6027), .Q(
        spi_master_clk_divider1[2]) );
  dfnrq1 \spi_master_clk_divider1_reg[1]  ( .D(N5644), .CP(n6042), .Q(
        spi_master_clk_divider1[1]) );
  dfnrq1 \spi_master_clk_divider1_reg[0]  ( .D(N5643), .CP(n6027), .Q(
        spi_master_clk_divider1[0]) );
  dfnrq1 multiregimpl1_regs0_reg ( .D(dbg_uart_dbg_uart_rx), .CP(n6075), .Q(
        multiregimpl1_regs0) );
  dfnrq1 multiregimpl1_regs1_reg ( .D(multiregimpl1_regs0), .CP(n6022), .Q(
        dbg_uart_rx_rx) );
  dfnrq1 multiregimpl0_regs0_reg ( .D(sys_uart_rx), .CP(n6055), .Q(
        multiregimpl0_regs0) );
  dfnrq1 multiregimpl0_regs1_reg ( .D(multiregimpl0_regs0), .CP(n6053), .Q(
        uart_phy_rx_rx) );
  dfnrq1 uart_phy_rx_rx_d_reg ( .D(N5704), .CP(n6051), .Q(uart_phy_rx_rx_d) );
  dfnrq1 rs232phy_rs232phyrx_state_reg ( .D(n3869), .CP(n6098), .Q(
        rs232phy_rs232phyrx_state) );
  dfnrq1 \uart_phy_rx_phase_reg[5]  ( .D(N3644), .CP(n6055), .Q(
        uart_phy_rx_phase[5]) );
  dfnrq1 \uart_phy_rx_phase_reg[6]  ( .D(N3645), .CP(n6053), .Q(
        uart_phy_rx_phase[6]) );
  dfnrq1 \uart_phy_rx_phase_reg[7]  ( .D(N3646), .CP(n6052), .Q(
        uart_phy_rx_phase[7]) );
  dfnrq1 \uart_phy_rx_phase_reg[8]  ( .D(N3647), .CP(n6052), .Q(
        uart_phy_rx_phase[8]) );
  dfnrq1 \uart_phy_rx_phase_reg[9]  ( .D(N3648), .CP(n6052), .Q(
        uart_phy_rx_phase[9]) );
  dfnrq1 \uart_phy_rx_phase_reg[10]  ( .D(N3649), .CP(n6052), .Q(
        uart_phy_rx_phase[10]) );
  dfnrq1 \uart_phy_rx_phase_reg[11]  ( .D(N3650), .CP(n6052), .Q(
        uart_phy_rx_phase[11]) );
  dfnrq1 \uart_phy_rx_phase_reg[12]  ( .D(N3651), .CP(n6052), .Q(
        uart_phy_rx_phase[12]) );
  dfnrq1 \uart_phy_rx_phase_reg[13]  ( .D(N3652), .CP(n6052), .Q(
        uart_phy_rx_phase[13]) );
  dfnrq1 \uart_phy_rx_phase_reg[14]  ( .D(N3653), .CP(n6052), .Q(
        uart_phy_rx_phase[14]) );
  dfnrq1 \uart_phy_rx_phase_reg[15]  ( .D(N3654), .CP(n6053), .Q(
        uart_phy_rx_phase[15]) );
  dfnrq1 \uart_phy_rx_phase_reg[16]  ( .D(N3655), .CP(n6022), .Q(
        uart_phy_rx_phase[16]) );
  dfnrq1 \uart_phy_rx_phase_reg[17]  ( .D(N3656), .CP(n6052), .Q(
        uart_phy_rx_phase[17]) );
  dfnrq1 \uart_phy_rx_phase_reg[18]  ( .D(N3657), .CP(n6075), .Q(
        uart_phy_rx_phase[18]) );
  dfnrq1 \uart_phy_rx_phase_reg[19]  ( .D(N3658), .CP(n6051), .Q(
        uart_phy_rx_phase[19]) );
  dfnrq1 \uart_phy_rx_phase_reg[20]  ( .D(N3659), .CP(n6075), .Q(
        uart_phy_rx_phase[20]) );
  dfnrq1 \uart_phy_rx_phase_reg[21]  ( .D(N3660), .CP(n6055), .Q(
        uart_phy_rx_phase[21]) );
  dfnrq1 \uart_phy_rx_phase_reg[22]  ( .D(N3661), .CP(n6053), .Q(
        uart_phy_rx_phase[22]) );
  dfnrq1 \uart_phy_rx_phase_reg[23]  ( .D(N3662), .CP(n6075), .Q(
        uart_phy_rx_phase[23]) );
  dfnrq1 \uart_phy_rx_phase_reg[24]  ( .D(N3663), .CP(n6053), .Q(
        uart_phy_rx_phase[24]) );
  dfnrq1 \uart_phy_rx_phase_reg[25]  ( .D(N3664), .CP(n6055), .Q(
        uart_phy_rx_phase[25]) );
  dfnrq1 \uart_phy_rx_phase_reg[26]  ( .D(N3665), .CP(n6053), .Q(
        uart_phy_rx_phase[26]) );
  dfnrq1 \uart_phy_rx_phase_reg[27]  ( .D(N3666), .CP(n6032), .Q(
        uart_phy_rx_phase[27]) );
  dfnrq1 \uart_phy_rx_phase_reg[28]  ( .D(N3667), .CP(n6051), .Q(
        uart_phy_rx_phase[28]) );
  dfnrq1 \uart_phy_rx_phase_reg[29]  ( .D(N3668), .CP(n6098), .Q(
        uart_phy_rx_phase[29]) );
  dfnrq1 \uart_phy_rx_phase_reg[30]  ( .D(N3669), .CP(n6075), .Q(
        uart_phy_rx_phase[30]) );
  dfnrq1 \uart_phy_rx_phase_reg[31]  ( .D(N3670), .CP(n6053), .Q(
        uart_phy_rx_phase[31]) );
  dfnrq1 uart_phy_rx_tick_reg ( .D(N5703), .CP(n6053), .Q(uart_phy_rx_tick) );
  dfnrq1 \uart_phy_rx_count_reg[0]  ( .D(n3868), .CP(n6053), .Q(
        uart_phy_rx_count[0]) );
  dfnrq1 \uart_phy_rx_count_reg[1]  ( .D(n3867), .CP(n6053), .Q(
        uart_phy_rx_count[1]) );
  dfnrq1 \uart_phy_rx_count_reg[2]  ( .D(n3866), .CP(n6053), .Q(
        uart_phy_rx_count[2]) );
  dfnrq1 \uart_phy_rx_count_reg[3]  ( .D(n3865), .CP(n6053), .Q(
        uart_phy_rx_count[3]) );
  dfnrq1 \uart_phy_rx_data_reg[7]  ( .D(n3722), .CP(n6053), .Q(
        uart_phy_rx_data[7]) );
  dfnrq1 \uart_phy_rx_data_reg[6]  ( .D(n3723), .CP(n6022), .Q(
        uart_phy_rx_data[6]) );
  dfnrq1 \uart_phy_rx_data_reg[5]  ( .D(n3724), .CP(n6032), .Q(
        uart_phy_rx_data[5]) );
  dfnrq1 \uart_phy_rx_data_reg[4]  ( .D(n3725), .CP(n6055), .Q(
        uart_phy_rx_data[4]) );
  dfnrq1 \uart_phy_rx_data_reg[3]  ( .D(n3726), .CP(n6053), .Q(
        uart_phy_rx_data[3]) );
  dfnrq1 \uart_phy_rx_data_reg[2]  ( .D(n3727), .CP(n6051), .Q(
        uart_phy_rx_data[2]) );
  dfnrq1 \uart_phy_rx_data_reg[1]  ( .D(n3728), .CP(n6022), .Q(
        uart_phy_rx_data[1]) );
  dfnrq1 \uart_phy_rx_data_reg[0]  ( .D(n3729), .CP(n6055), .Q(
        uart_phy_rx_data[0]) );
  dfnrq1 dbg_uart_rx_rx_d_reg ( .D(N5758), .CP(n6055), .Q(dbg_uart_rx_rx_d) );
  dfnrq1 multiregimpl2_regs0_reg ( .D(gpio_in_pad), .CP(n6098), .Q(
        multiregimpl2_regs0) );
  dfnrq1 multiregimpl2_regs1_reg ( .D(multiregimpl2_regs0), .CP(n6023), .Q(
        csrbank5_in_w) );
  dfnrq1 \dbg_uart_rx_count_reg[0]  ( .D(n3881), .CP(n6058), .Q(
        dbg_uart_rx_count[0]) );
  dfnrq1 uartwishbonebridge_rs232phyrx_state_reg ( .D(n3882), .CP(n6098), .Q(
        uartwishbonebridge_rs232phyrx_state) );
  dfnrq1 dbg_uart_rx_tick_reg ( .D(N5757), .CP(n6116), .Q(dbg_uart_rx_tick) );
  dfnrq1 \dbg_uart_rx_phase_reg[0]  ( .D(N5046), .CP(n6115), .Q(
        dbg_uart_rx_phase[0]) );
  dfnrq1 \dbg_uart_rx_phase_reg[1]  ( .D(N5047), .CP(n6116), .Q(
        dbg_uart_rx_phase[1]) );
  dfnrq1 \dbg_uart_rx_phase_reg[2]  ( .D(N5048), .CP(n6116), .Q(
        dbg_uart_rx_phase[2]) );
  dfnrq1 \dbg_uart_rx_phase_reg[3]  ( .D(N5049), .CP(n6116), .Q(
        dbg_uart_rx_phase[3]) );
  dfnrq1 \dbg_uart_rx_phase_reg[4]  ( .D(N5050), .CP(n6062), .Q(
        dbg_uart_rx_phase[4]) );
  dfnrq1 \dbg_uart_rx_phase_reg[5]  ( .D(N5051), .CP(n6022), .Q(
        dbg_uart_rx_phase[5]) );
  dfnrq1 \dbg_uart_rx_phase_reg[6]  ( .D(N5052), .CP(n6116), .Q(
        dbg_uart_rx_phase[6]) );
  dfnrq1 \dbg_uart_rx_phase_reg[7]  ( .D(N5053), .CP(n6045), .Q(
        dbg_uart_rx_phase[7]) );
  dfnrq1 \dbg_uart_rx_phase_reg[8]  ( .D(N5054), .CP(n6115), .Q(
        dbg_uart_rx_phase[8]) );
  dfnrq1 \dbg_uart_rx_phase_reg[9]  ( .D(N5055), .CP(n6044), .Q(
        dbg_uart_rx_phase[9]) );
  dfnrq1 \dbg_uart_rx_phase_reg[10]  ( .D(N5056), .CP(n6116), .Q(
        dbg_uart_rx_phase[10]) );
  dfnrq1 \dbg_uart_rx_phase_reg[11]  ( .D(N5057), .CP(n6023), .Q(
        dbg_uart_rx_phase[11]) );
  dfnrq1 \dbg_uart_rx_phase_reg[12]  ( .D(N5058), .CP(n6116), .Q(
        dbg_uart_rx_phase[12]) );
  dfnrq1 \dbg_uart_rx_phase_reg[13]  ( .D(N5059), .CP(n6032), .Q(
        dbg_uart_rx_phase[13]) );
  dfnrq1 \dbg_uart_rx_phase_reg[14]  ( .D(N5060), .CP(n6116), .Q(
        dbg_uart_rx_phase[14]) );
  dfnrq1 \dbg_uart_rx_phase_reg[15]  ( .D(N5061), .CP(n6115), .Q(
        dbg_uart_rx_phase[15]) );
  dfnrq1 \dbg_uart_rx_phase_reg[16]  ( .D(N5062), .CP(n6128), .Q(
        dbg_uart_rx_phase[16]) );
  dfnrq1 \dbg_uart_rx_phase_reg[17]  ( .D(N5063), .CP(n6115), .Q(
        dbg_uart_rx_phase[17]) );
  dfnrq1 \dbg_uart_rx_phase_reg[18]  ( .D(N5064), .CP(n6116), .Q(
        dbg_uart_rx_phase[18]) );
  dfnrq1 \dbg_uart_rx_phase_reg[19]  ( .D(N5065), .CP(n6116), .Q(
        dbg_uart_rx_phase[19]) );
  dfnrq1 \dbg_uart_rx_phase_reg[20]  ( .D(N5066), .CP(n6098), .Q(
        dbg_uart_rx_phase[20]) );
  dfnrq1 \dbg_uart_rx_phase_reg[21]  ( .D(N5067), .CP(n6026), .Q(
        dbg_uart_rx_phase[21]) );
  dfnrq1 \dbg_uart_rx_phase_reg[22]  ( .D(N5068), .CP(n6115), .Q(
        dbg_uart_rx_phase[22]) );
  dfnrq1 \dbg_uart_rx_phase_reg[23]  ( .D(N5069), .CP(n6051), .Q(
        dbg_uart_rx_phase[23]) );
  dfnrq1 \dbg_uart_rx_phase_reg[24]  ( .D(N5070), .CP(n6054), .Q(
        dbg_uart_rx_phase[24]) );
  dfnrq1 \dbg_uart_rx_phase_reg[25]  ( .D(N5071), .CP(n6029), .Q(
        dbg_uart_rx_phase[25]) );
  dfnrq1 \dbg_uart_rx_phase_reg[26]  ( .D(N5072), .CP(n6116), .Q(
        dbg_uart_rx_phase[26]) );
  dfnrq1 \dbg_uart_rx_phase_reg[27]  ( .D(N5073), .CP(n6059), .Q(
        dbg_uart_rx_phase[27]) );
  dfnrq1 \dbg_uart_rx_phase_reg[28]  ( .D(N5074), .CP(n6060), .Q(
        dbg_uart_rx_phase[28]) );
  dfnrq1 \dbg_uart_rx_phase_reg[29]  ( .D(N5075), .CP(n6061), .Q(
        dbg_uart_rx_phase[29]) );
  dfnrq1 \dbg_uart_rx_phase_reg[30]  ( .D(N5076), .CP(n6062), .Q(
        dbg_uart_rx_phase[30]) );
  dfnrq1 \dbg_uart_rx_phase_reg[31]  ( .D(N5077), .CP(n6056), .Q(
        dbg_uart_rx_phase[31]) );
  dfnrq1 \dbg_uart_rx_count_reg[1]  ( .D(n3880), .CP(n6054), .Q(
        dbg_uart_rx_count[1]) );
  dfnrq1 \dbg_uart_rx_count_reg[2]  ( .D(n3879), .CP(n6061), .Q(
        dbg_uart_rx_count[2]) );
  dfnrq1 \dbg_uart_rx_count_reg[3]  ( .D(n3878), .CP(n6059), .Q(
        dbg_uart_rx_count[3]) );
  dfnrq1 \dbg_uart_rx_data_reg[7]  ( .D(n3870), .CP(n6062), .Q(
        dbg_uart_rx_data[7]) );
  dfnrq1 \dbg_uart_rx_data_reg[6]  ( .D(n3871), .CP(n6056), .Q(
        dbg_uart_rx_data[6]) );
  dfnrq1 \dbg_uart_rx_data_reg[5]  ( .D(n3872), .CP(n6054), .Q(
        dbg_uart_rx_data[5]) );
  dfnrq1 \dbg_uart_rx_data_reg[4]  ( .D(n3873), .CP(n6060), .Q(
        dbg_uart_rx_data[4]) );
  dfnrq1 \dbg_uart_rx_data_reg[3]  ( .D(n3874), .CP(n6056), .Q(
        dbg_uart_rx_data[3]) );
  dfnrq1 \dbg_uart_rx_data_reg[2]  ( .D(n3875), .CP(n6060), .Q(
        dbg_uart_rx_data[2]) );
  dfnrq1 \dbg_uart_rx_data_reg[1]  ( .D(n3876), .CP(n6058), .Q(
        dbg_uart_rx_data[1]) );
  dfnrq1 \dbg_uart_rx_data_reg[0]  ( .D(n3877), .CP(n6062), .Q(
        dbg_uart_rx_data[0]) );
  dfnrq1 gpioin3_gpioin3_in_pads_n_d_reg ( .D(N6228), .CP(n6056), .Q(
        gpioin3_gpioin3_in_pads_n_d) );
  dfnrq1 gpioin4_gpioin4_in_pads_n_d_reg ( .D(N6236), .CP(n6061), .Q(
        gpioin4_gpioin4_in_pads_n_d) );
  dfnrq1 gpioin5_gpioin5_in_pads_n_d_reg ( .D(N6244), .CP(n6062), .Q(
        gpioin5_gpioin5_in_pads_n_d) );
  dfnrq1 \memdat_3_reg[0]  ( .D(n4546), .CP(n6047), .Q(
        uart_rx_fifo_fifo_out_payload_data[0]) );
  dfnrq1 \interface11_bank_bus_dat_r_reg[0]  ( .D(N4772), .CP(n6037), .Q(
        interface11_bank_bus_dat_r[0]) );
  dfnrq1 \dbg_uart_data_reg[0]  ( .D(n3283), .CP(n6038), .Q(
        dbg_uart_wishbone_dat_w[0]) );
  dfnrq1 \dbg_uart_data_reg[8]  ( .D(n3275), .CP(n6048), .Q(
        dbg_uart_wishbone_dat_w[8]) );
  dfnrq1 \dbg_uart_data_reg[16]  ( .D(n3267), .CP(n6038), .Q(
        dbg_uart_wishbone_dat_w[16]) );
  dfnrq1 \dbg_uart_data_reg[24]  ( .D(n3259), .CP(n6039), .Q(
        dbg_uart_wishbone_dat_w[24]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[24]  ( .D(n3303), .CP(n6048), .Q(
        csrbank0_scratch0_w[24]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[24]  ( .D(N4123), .CP(n6036), .Q(
        interface0_bank_bus_dat_r[24]) );
  dfnrq1 mgmtsoc_vexriscv_reset_debug_logic_reg ( .D(N5281), .CP(n6041), .Q(
        mgmtsoc_vexriscv_reset_debug_logic) );
  dfnrq1 mgmtsoc_vexriscv_debug_reset_reg ( .D(N5235), .CP(n6036), .Q(
        mgmtsoc_vexriscv_debug_reset) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[0]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[0]), .CP(n6038), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[0]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[1]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[1]), .CP(n6037), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[1]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[2]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[2]), .CP(n6037), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[2]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[3]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[3]), .CP(n6114), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[3]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[4]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[4]), .CP(n6047), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[4]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[5]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[5]), .CP(n6114), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[5]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[6]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[6]), .CP(n6114), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[6]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[7]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[7]), .CP(n6114), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[7]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[8]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[8]), .CP(n6037), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[8]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[9]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[9]), .CP(n6114), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[9]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[10]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[10]), .CP(n6114), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[10]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[11]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[11]), .CP(n6037), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[11]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[12]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[12]), .CP(n6047), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[12]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[13]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[13]), .CP(n6038), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[13]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[14]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[14]), .CP(n6039), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[14]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[15]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[15]), .CP(n6048), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[15]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[16]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[16]), .CP(n6036), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[16]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[17]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[17]), .CP(n6041), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[17]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[18]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[18]), .CP(n6044), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[18]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[19]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[19]), .CP(n6044), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[19]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[20]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[20]), .CP(n6044), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[20]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[21]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[21]), .CP(n6044), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[21]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[22]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[22]), .CP(n6044), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[22]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[23]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[23]), .CP(n6044), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[23]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[24]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[24]), .CP(n6044), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[24]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[25]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[25]), .CP(n6044), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[25]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[26]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[26]), .CP(n6045), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[26]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[27]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[27]), .CP(n6045), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[27]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[28]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[28]), .CP(n6045), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[28]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[29]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[29]), .CP(n6045), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[29]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[30]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[30]), .CP(n6045), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[30]) );
  dfnrq1 \mgmtsoc_vexriscv_debug_bus_dat_r_reg[31]  ( .D(
        mgmtsoc_vexriscv_o_rsp_data[31]), .CP(n6045), .Q(
        mgmtsoc_vexriscv_debug_bus_dat_r[31]) );
  dfnrq1 mgmtsoc_vexriscv_i_cmd_valid_reg ( .D(n3360), .CP(n6045), .Q(
        mgmtsoc_vexriscv_i_cmd_valid) );
  dfnrq1 mgmtsoc_vexriscv_transfer_complete_reg ( .D(n3400), .CP(n6045), .Q(
        mgmtsoc_vexriscv_transfer_complete) );
  dfnrq1 mgmtsoc_vexriscv_debug_bus_ack_reg ( .D(n3402), .CP(n6046), .Q(
        mgmtsoc_vexriscv_debug_bus_ack) );
  dfnrq1 \uartwishbonebridge_state_reg[0]  ( .D(N6262), .CP(n6046), .Q(
        uartwishbonebridge_state[0]) );
  dfnrq1 uartwishbonebridge_rs232phytx_state_reg ( .D(n3097), .CP(n6046), .Q(
        uartwishbonebridge_rs232phytx_state) );
  dfnrq1 \dbg_uart_tx_phase_reg[0]  ( .D(N5014), .CP(n6046), .Q(
        dbg_uart_tx_phase[0]) );
  dfnrq1 \dbg_uart_tx_phase_reg[1]  ( .D(N5015), .CP(n6046), .Q(
        dbg_uart_tx_phase[1]) );
  dfnrq1 \dbg_uart_tx_phase_reg[2]  ( .D(N5016), .CP(n6046), .Q(
        dbg_uart_tx_phase[2]) );
  dfnrq1 \dbg_uart_tx_phase_reg[7]  ( .D(N5021), .CP(n6046), .Q(
        dbg_uart_tx_phase[7]) );
  dfnrq1 \dbg_uart_tx_phase_reg[8]  ( .D(N5022), .CP(n6046), .Q(
        dbg_uart_tx_phase[8]) );
  dfnrq1 \dbg_uart_tx_phase_reg[11]  ( .D(N5025), .CP(n6047), .Q(
        dbg_uart_tx_phase[11]) );
  dfnrq1 \dbg_uart_tx_phase_reg[12]  ( .D(N5026), .CP(n6047), .Q(
        dbg_uart_tx_phase[12]) );
  dfnrq1 \dbg_uart_tx_phase_reg[13]  ( .D(N5027), .CP(n6047), .Q(
        dbg_uart_tx_phase[13]) );
  dfnrq1 \dbg_uart_tx_phase_reg[14]  ( .D(N5028), .CP(n6047), .Q(
        dbg_uart_tx_phase[14]) );
  dfnrq1 \dbg_uart_tx_phase_reg[15]  ( .D(N5029), .CP(n6047), .Q(
        dbg_uart_tx_phase[15]) );
  dfnrq1 \dbg_uart_tx_phase_reg[17]  ( .D(N5031), .CP(n6047), .Q(
        dbg_uart_tx_phase[17]) );
  dfnrq1 \dbg_uart_tx_phase_reg[20]  ( .D(N5034), .CP(n6047), .Q(
        dbg_uart_tx_phase[20]) );
  dfnrq1 \dbg_uart_tx_phase_reg[21]  ( .D(N5035), .CP(n6094), .Q(
        dbg_uart_tx_phase[21]) );
  dfnrq1 \dbg_uart_tx_phase_reg[22]  ( .D(N5036), .CP(n6047), .Q(
        dbg_uart_tx_phase[22]) );
  dfnrq1 \dbg_uart_tx_phase_reg[23]  ( .D(N5037), .CP(n6114), .Q(
        dbg_uart_tx_phase[23]) );
  dfnrq1 \dbg_uart_tx_phase_reg[25]  ( .D(N5039), .CP(n6057), .Q(
        dbg_uart_tx_phase[25]) );
  dfnrq1 dbg_uart_tx_tick_reg ( .D(N5756), .CP(n6113), .Q(dbg_uart_tx_tick) );
  dfnrq1 \dbg_uart_tx_phase_reg[3]  ( .D(N5017), .CP(n6094), .Q(
        dbg_uart_tx_phase[3]) );
  dfnrq1 \dbg_uart_tx_phase_reg[4]  ( .D(N5018), .CP(n6095), .Q(
        dbg_uart_tx_phase[4]) );
  dfnrq1 \dbg_uart_tx_phase_reg[5]  ( .D(N5019), .CP(n6102), .Q(
        dbg_uart_tx_phase[5]) );
  dfnrq1 \dbg_uart_tx_phase_reg[6]  ( .D(N5020), .CP(n6048), .Q(
        dbg_uart_tx_phase[6]) );
  dfnrq1 \dbg_uart_tx_phase_reg[9]  ( .D(N5023), .CP(n6048), .Q(
        dbg_uart_tx_phase[9]) );
  dfnrq1 \dbg_uart_tx_phase_reg[10]  ( .D(N5024), .CP(n6048), .Q(
        dbg_uart_tx_phase[10]) );
  dfnrq1 \dbg_uart_tx_phase_reg[16]  ( .D(N5030), .CP(n6048), .Q(
        dbg_uart_tx_phase[16]) );
  dfnrq1 \dbg_uart_tx_phase_reg[18]  ( .D(N5032), .CP(n6048), .Q(
        dbg_uart_tx_phase[18]) );
  dfnrq1 \dbg_uart_tx_phase_reg[19]  ( .D(N5033), .CP(n6048), .Q(
        dbg_uart_tx_phase[19]) );
  dfnrq1 \dbg_uart_tx_phase_reg[24]  ( .D(N5038), .CP(n6048), .Q(
        dbg_uart_tx_phase[24]) );
  dfnrq1 \dbg_uart_tx_phase_reg[26]  ( .D(N5040), .CP(n6048), .Q(
        dbg_uart_tx_phase[26]) );
  dfnrq1 \dbg_uart_tx_phase_reg[27]  ( .D(N5041), .CP(n6049), .Q(
        dbg_uart_tx_phase[27]) );
  dfnrq1 \dbg_uart_tx_phase_reg[28]  ( .D(N5042), .CP(n6049), .Q(
        dbg_uart_tx_phase[28]) );
  dfnrq1 \dbg_uart_tx_phase_reg[29]  ( .D(N5043), .CP(n6049), .Q(
        dbg_uart_tx_phase[29]) );
  dfnrq1 \dbg_uart_tx_phase_reg[30]  ( .D(N5044), .CP(n6049), .Q(
        dbg_uart_tx_phase[30]) );
  dfnrq1 \dbg_uart_tx_phase_reg[31]  ( .D(N5045), .CP(n6049), .Q(
        dbg_uart_tx_phase[31]) );
  dfnrq1 \dbg_uart_tx_count_reg[0]  ( .D(n3101), .CP(n6049), .Q(
        dbg_uart_tx_count[0]) );
  dfnrq1 \dbg_uart_tx_count_reg[1]  ( .D(n3100), .CP(n6049), .Q(
        dbg_uart_tx_count[1]) );
  dfnrq1 \dbg_uart_tx_count_reg[2]  ( .D(n3099), .CP(n6049), .Q(
        dbg_uart_tx_count[2]) );
  dfnrq1 \dbg_uart_tx_count_reg[3]  ( .D(n3098), .CP(n6038), .Q(
        dbg_uart_tx_count[3]) );
  dfnrq1 \uartwishbonebridge_state_reg[2]  ( .D(N6264), .CP(n6102), .Q(
        uartwishbonebridge_state[2]) );
  dfnrq1 \dbg_uart_count_reg[0]  ( .D(n4088), .CP(n6040), .Q(dbg_uart_count[0]) );
  dfnrq1 \dbg_uart_count_reg[15]  ( .D(n4083), .CP(n6113), .Q(
        dbg_uart_count[15]) );
  dfnrq1 \dbg_uart_count_reg[13]  ( .D(n4081), .CP(n6092), .Q(
        dbg_uart_count[13]) );
  dfnrq1 \dbg_uart_count_reg[12]  ( .D(n4080), .CP(n6041), .Q(
        dbg_uart_count[12]) );
  dfnrq1 \dbg_uart_count_reg[11]  ( .D(n4079), .CP(n6114), .Q(
        dbg_uart_count[11]) );
  dfnrq1 \dbg_uart_count_reg[10]  ( .D(n4078), .CP(n6102), .Q(
        dbg_uart_count[10]) );
  dfnrq1 \dbg_uart_count_reg[8]  ( .D(n4076), .CP(n6050), .Q(dbg_uart_count[8]) );
  dfnrq1 \dbg_uart_count_reg[7]  ( .D(n4075), .CP(n6052), .Q(dbg_uart_count[7]) );
  dfnrq1 \dbg_uart_count_reg[5]  ( .D(n4073), .CP(n6050), .Q(dbg_uart_count[5]) );
  dfnrq1 \dbg_uart_count_reg[4]  ( .D(n4072), .CP(n6115), .Q(dbg_uart_count[4]) );
  dfnrq1 \dbg_uart_count_reg[3]  ( .D(n4071), .CP(n6115), .Q(dbg_uart_count[3]) );
  dfnrq1 \dbg_uart_count_reg[2]  ( .D(n4070), .CP(n6115), .Q(dbg_uart_count[2]) );
  dfnrq1 \dbg_uart_count_reg[1]  ( .D(n4069), .CP(n6052), .Q(dbg_uart_count[1]) );
  dfnrq1 \dbg_uart_count_reg[19]  ( .D(n4087), .CP(n6050), .Q(
        dbg_uart_count[19]) );
  dfnrq1 \dbg_uart_count_reg[18]  ( .D(n4086), .CP(n6115), .Q(
        dbg_uart_count[18]) );
  dfnrq1 \dbg_uart_count_reg[17]  ( .D(n4085), .CP(n6115), .Q(
        dbg_uart_count[17]) );
  dfnrq1 \dbg_uart_count_reg[16]  ( .D(n4084), .CP(n6052), .Q(
        dbg_uart_count[16]) );
  dfnrq1 \dbg_uart_count_reg[14]  ( .D(n4082), .CP(n6050), .Q(
        dbg_uart_count[14]) );
  dfnrq1 \dbg_uart_count_reg[9]  ( .D(n4077), .CP(n6115), .Q(dbg_uart_count[9]) );
  dfnrq1 \dbg_uart_count_reg[6]  ( .D(n4074), .CP(n6052), .Q(dbg_uart_count[6]) );
  dfnrq1 \dbg_uart_cmd_reg[0]  ( .D(n3117), .CP(n6052), .Q(dbg_uart_cmd[0]) );
  dfnrq1 \dbg_uart_cmd_reg[1]  ( .D(n3116), .CP(n6050), .Q(dbg_uart_cmd[1]) );
  dfnrq1 \dbg_uart_cmd_reg[2]  ( .D(n3115), .CP(n6115), .Q(dbg_uart_cmd[2]) );
  dfnrq1 \dbg_uart_cmd_reg[3]  ( .D(n3114), .CP(n6052), .Q(dbg_uart_cmd[3]) );
  dfnrq1 \dbg_uart_cmd_reg[4]  ( .D(n3113), .CP(n6050), .Q(dbg_uart_cmd[4]) );
  dfnrq1 \dbg_uart_cmd_reg[5]  ( .D(n3112), .CP(n6115), .Q(dbg_uart_cmd[5]) );
  dfnrq1 \dbg_uart_cmd_reg[6]  ( .D(n3111), .CP(n6052), .Q(dbg_uart_cmd[6]) );
  dfnrq1 \dbg_uart_cmd_reg[7]  ( .D(n3110), .CP(n6050), .Q(dbg_uart_cmd[7]) );
  dfnrq1 \uartwishbonebridge_state_reg[1]  ( .D(N6263), .CP(n6115), .Q(
        uartwishbonebridge_state[1]) );
  dfnrq1 \dbg_uart_bytes_count_reg[0]  ( .D(n3285), .CP(n6052), .Q(
        dbg_uart_bytes_count[0]) );
  dfnrq1 \dbg_uart_bytes_count_reg[1]  ( .D(n3284), .CP(n6050), .Q(
        dbg_uart_bytes_count[1]) );
  dfnrq1 \grant_reg[1]  ( .D(n4516), .CP(n6050), .Q(grant[1]) );
  dfnrq1 \grant_reg[0]  ( .D(n4517), .CP(n6050), .Q(grant[0]) );
  dfnrq1 \count_reg[0]  ( .D(n4537), .CP(n6050), .Q(count[0]) );
  dfnrq1 \count_reg[19]  ( .D(n4536), .CP(n6063), .Q(count[19]) );
  dfnrq1 \count_reg[18]  ( .D(n4535), .CP(n6060), .Q(count[18]) );
  dfnrq1 \count_reg[17]  ( .D(n4534), .CP(n6060), .Q(count[17]) );
  dfnrq1 \count_reg[16]  ( .D(n4533), .CP(n6060), .Q(count[16]) );
  dfnrq1 \count_reg[15]  ( .D(n4532), .CP(n6060), .Q(count[15]) );
  dfnrq1 \count_reg[14]  ( .D(n4531), .CP(n6060), .Q(count[14]) );
  dfnrq1 \count_reg[13]  ( .D(n4530), .CP(n6061), .Q(count[13]) );
  dfnrq1 \count_reg[12]  ( .D(n4529), .CP(n6061), .Q(count[12]) );
  dfnrq1 \count_reg[11]  ( .D(n4528), .CP(n6061), .Q(count[11]) );
  dfnrq1 \count_reg[10]  ( .D(n4527), .CP(n6061), .Q(count[10]) );
  dfnrq1 \count_reg[9]  ( .D(n4526), .CP(n6061), .Q(count[9]) );
  dfnrq1 \count_reg[8]  ( .D(n4525), .CP(n6061), .Q(count[8]) );
  dfnrq1 \count_reg[7]  ( .D(n4524), .CP(n6061), .Q(count[7]) );
  dfnrq1 \count_reg[6]  ( .D(n4523), .CP(n6061), .Q(count[6]) );
  dfnrq1 \count_reg[5]  ( .D(n4522), .CP(n6062), .Q(count[5]) );
  dfnrq1 \count_reg[4]  ( .D(n4521), .CP(n6062), .Q(count[4]) );
  dfnrq1 \count_reg[3]  ( .D(n4520), .CP(n6062), .Q(count[3]) );
  dfnrq1 \count_reg[2]  ( .D(n4519), .CP(n6062), .Q(count[2]) );
  dfnrq1 \count_reg[1]  ( .D(n4518), .CP(n6062), .Q(count[1]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[0]  ( .D(n3359), .CP(n6062), .Q(
        mgmtsoc_bus_errors_status[0]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[31]  ( .D(n3358), .CP(n6062), .Q(
        mgmtsoc_bus_errors_status[31]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[30]  ( .D(n3357), .CP(n6062), .Q(
        mgmtsoc_bus_errors_status[30]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[29]  ( .D(n3356), .CP(n6028), .Q(
        mgmtsoc_bus_errors_status[29]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[28]  ( .D(n3355), .CP(n6099), .Q(
        mgmtsoc_bus_errors_status[28]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[27]  ( .D(n3354), .CP(n6028), .Q(
        mgmtsoc_bus_errors_status[27]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[26]  ( .D(n3353), .CP(n6099), .Q(
        mgmtsoc_bus_errors_status[26]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[25]  ( .D(n3352), .CP(n6028), .Q(
        mgmtsoc_bus_errors_status[25]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[24]  ( .D(n3351), .CP(n6099), .Q(
        mgmtsoc_bus_errors_status[24]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[23]  ( .D(n3350), .CP(n6028), .Q(
        mgmtsoc_bus_errors_status[23]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[22]  ( .D(n3349), .CP(n6099), .Q(
        mgmtsoc_bus_errors_status[22]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[21]  ( .D(n3348), .CP(n6063), .Q(
        mgmtsoc_bus_errors_status[21]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[20]  ( .D(n3347), .CP(n6063), .Q(
        mgmtsoc_bus_errors_status[20]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[19]  ( .D(n3346), .CP(n6118), .Q(
        mgmtsoc_bus_errors_status[19]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[18]  ( .D(n3345), .CP(n6073), .Q(
        mgmtsoc_bus_errors_status[18]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[17]  ( .D(n3344), .CP(n6063), .Q(
        mgmtsoc_bus_errors_status[17]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[16]  ( .D(n3343), .CP(n6118), .Q(
        mgmtsoc_bus_errors_status[16]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[15]  ( .D(n3342), .CP(n6063), .Q(
        mgmtsoc_bus_errors_status[15]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[14]  ( .D(n3341), .CP(n6065), .Q(
        mgmtsoc_bus_errors_status[14]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[13]  ( .D(n3340), .CP(n6023), .Q(
        mgmtsoc_bus_errors_status[13]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[12]  ( .D(n3339), .CP(n6117), .Q(
        mgmtsoc_bus_errors_status[12]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[11]  ( .D(n3338), .CP(n6118), .Q(
        mgmtsoc_bus_errors_status[11]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[10]  ( .D(n3337), .CP(n6120), .Q(
        mgmtsoc_bus_errors_status[10]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[9]  ( .D(n3336), .CP(n6063), .Q(
        mgmtsoc_bus_errors_status[9]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[8]  ( .D(n3335), .CP(n6065), .Q(
        mgmtsoc_bus_errors_status[8]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[7]  ( .D(n3334), .CP(n6064), .Q(
        mgmtsoc_bus_errors_status[7]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[6]  ( .D(n3333), .CP(n6070), .Q(
        mgmtsoc_bus_errors_status[6]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[5]  ( .D(n3332), .CP(n6040), .Q(
        mgmtsoc_bus_errors_status[5]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[4]  ( .D(n3331), .CP(n6027), .Q(
        mgmtsoc_bus_errors_status[4]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[3]  ( .D(n3330), .CP(n6027), .Q(
        mgmtsoc_bus_errors_status[3]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[2]  ( .D(n3329), .CP(n6113), .Q(
        mgmtsoc_bus_errors_status[2]) );
  dfnrq1 \mgmtsoc_bus_errors_reg[1]  ( .D(n3328), .CP(n6113), .Q(
        mgmtsoc_bus_errors_status[1]) );
  dfnrq1 dbg_uart_incr_reg ( .D(n4068), .CP(n6027), .Q(dbg_uart_incr) );
  dfnrq1 \dbg_uart_length_reg[0]  ( .D(n3109), .CP(n6113), .Q(
        dbg_uart_length[0]) );
  dfnrq1 \dbg_uart_length_reg[1]  ( .D(n3108), .CP(n6027), .Q(
        dbg_uart_length[1]) );
  dfnrq1 \dbg_uart_length_reg[2]  ( .D(n3107), .CP(n6063), .Q(
        dbg_uart_length[2]) );
  dfnrq1 \dbg_uart_length_reg[3]  ( .D(n3106), .CP(n6063), .Q(
        dbg_uart_length[3]) );
  dfnrq1 \dbg_uart_length_reg[4]  ( .D(n3105), .CP(n6063), .Q(
        dbg_uart_length[4]) );
  dfnrq1 \dbg_uart_length_reg[5]  ( .D(n3104), .CP(n6063), .Q(
        dbg_uart_length[5]) );
  dfnrq1 \dbg_uart_length_reg[6]  ( .D(n3103), .CP(n6063), .Q(
        dbg_uart_length[6]) );
  dfnrq1 \dbg_uart_length_reg[7]  ( .D(n3102), .CP(n6063), .Q(
        dbg_uart_length[7]) );
  dfnrq1 \dbg_uart_words_count_reg[0]  ( .D(n3293), .CP(n6063), .Q(
        dbg_uart_words_count[0]) );
  dfnrq1 \dbg_uart_words_count_reg[1]  ( .D(n3292), .CP(n6064), .Q(
        dbg_uart_words_count[1]) );
  dfnrq1 \dbg_uart_words_count_reg[2]  ( .D(n3291), .CP(n6064), .Q(
        dbg_uart_words_count[2]) );
  dfnrq1 \dbg_uart_words_count_reg[3]  ( .D(n3290), .CP(n6064), .Q(
        dbg_uart_words_count[3]) );
  dfnrq1 \dbg_uart_words_count_reg[4]  ( .D(n3289), .CP(n6064), .Q(
        dbg_uart_words_count[4]) );
  dfnrq1 \dbg_uart_words_count_reg[5]  ( .D(n3288), .CP(n6064), .Q(
        dbg_uart_words_count[5]) );
  dfnrq1 \dbg_uart_words_count_reg[6]  ( .D(n3287), .CP(n6064), .Q(
        dbg_uart_words_count[6]) );
  dfnrq1 \dbg_uart_words_count_reg[7]  ( .D(n3286), .CP(n6064), .Q(
        dbg_uart_words_count[7]) );
  dfnrq1 \dbg_uart_address_reg[0]  ( .D(n3251), .CP(n6064), .Q(
        dbg_uart_wishbone_adr[0]) );
  dfnrq1 \dbg_uart_address_reg[1]  ( .D(n3250), .CP(n6063), .Q(
        dbg_uart_wishbone_adr[1]) );
  dfnrq1 \dbg_uart_address_reg[2]  ( .D(n3249), .CP(n6118), .Q(
        dbg_uart_wishbone_adr[2]) );
  dfnrq1 \dbg_uart_address_reg[3]  ( .D(n3248), .CP(n6118), .Q(
        dbg_uart_wishbone_adr[3]) );
  dfnrq1 \dbg_uart_address_reg[4]  ( .D(n3247), .CP(n6063), .Q(
        dbg_uart_wishbone_adr[4]) );
  dfnrq1 \dbg_uart_address_reg[5]  ( .D(n3246), .CP(n6070), .Q(
        dbg_uart_wishbone_adr[5]) );
  dfnrq1 \dbg_uart_address_reg[6]  ( .D(n3245), .CP(n6118), .Q(
        dbg_uart_wishbone_adr[6]) );
  dfnrq1 \dbg_uart_address_reg[7]  ( .D(n3244), .CP(n6063), .Q(
        dbg_uart_wishbone_adr[7]) );
  dfnrq1 \dbg_uart_address_reg[8]  ( .D(n3243), .CP(n6064), .Q(
        dbg_uart_wishbone_adr[8]) );
  dfnrq1 \dbg_uart_address_reg[9]  ( .D(n3242), .CP(n6065), .Q(
        dbg_uart_wishbone_adr[9]) );
  dfnrq1 \dbg_uart_address_reg[10]  ( .D(n3241), .CP(n6065), .Q(
        dbg_uart_wishbone_adr[10]) );
  dfnrq1 \dbg_uart_address_reg[11]  ( .D(n3240), .CP(n6065), .Q(
        dbg_uart_wishbone_adr[11]) );
  dfnrq1 \dbg_uart_address_reg[12]  ( .D(n3239), .CP(n6065), .Q(
        dbg_uart_wishbone_adr[12]) );
  dfnrq1 \dbg_uart_address_reg[13]  ( .D(n3238), .CP(n6065), .Q(
        dbg_uart_wishbone_adr[13]) );
  dfnrq1 \dbg_uart_address_reg[14]  ( .D(n3237), .CP(n6065), .Q(
        dbg_uart_wishbone_adr[14]) );
  dfnrq1 \dbg_uart_address_reg[15]  ( .D(n3236), .CP(n6065), .Q(
        dbg_uart_wishbone_adr[15]) );
  dfnrq1 \dbg_uart_address_reg[16]  ( .D(n3235), .CP(n6065), .Q(
        dbg_uart_wishbone_adr[16]) );
  dfnrq1 \dbg_uart_address_reg[17]  ( .D(n3234), .CP(n6066), .Q(
        dbg_uart_wishbone_adr[17]) );
  dfnrq1 \dbg_uart_address_reg[18]  ( .D(n3233), .CP(n6066), .Q(
        dbg_uart_wishbone_adr[18]) );
  dfnrq1 \dbg_uart_address_reg[19]  ( .D(n3232), .CP(n6066), .Q(
        dbg_uart_wishbone_adr[19]) );
  dfnrq1 \dbg_uart_address_reg[20]  ( .D(n3231), .CP(n6066), .Q(
        dbg_uart_wishbone_adr[20]) );
  dfnrq1 \dbg_uart_address_reg[21]  ( .D(n3230), .CP(n6066), .Q(
        dbg_uart_wishbone_adr[21]) );
  dfnrq1 \dbg_uart_address_reg[22]  ( .D(n3229), .CP(n6066), .Q(
        dbg_uart_wishbone_adr[22]) );
  dfnrq1 \dbg_uart_address_reg[23]  ( .D(n3228), .CP(n6066), .Q(
        dbg_uart_wishbone_adr[23]) );
  dfnrq1 \dbg_uart_address_reg[24]  ( .D(n3227), .CP(n6066), .Q(
        dbg_uart_wishbone_adr[24]) );
  dfnrq1 \dbg_uart_address_reg[25]  ( .D(n3226), .CP(n6066), .Q(
        dbg_uart_wishbone_adr[25]) );
  dfnrq1 \dbg_uart_address_reg[26]  ( .D(n3225), .CP(n6120), .Q(
        dbg_uart_wishbone_adr[26]) );
  dfnrq1 \dbg_uart_address_reg[27]  ( .D(n3224), .CP(n6117), .Q(
        dbg_uart_wishbone_adr[27]) );
  dfnrq1 \dbg_uart_address_reg[28]  ( .D(n3223), .CP(n6117), .Q(
        dbg_uart_wishbone_adr[28]) );
  dfnrq1 \dbg_uart_address_reg[29]  ( .D(n3222), .CP(n6117), .Q(
        dbg_uart_wishbone_adr[29]) );
  dfnrq1 \slave_sel_r_reg[4]  ( .D(N6302), .CP(n6117), .Q(slave_sel_r[4]) );
  dfnrq1 \slave_sel_r_reg[2]  ( .D(N6300), .CP(n6068), .Q(slave_sel_r[2]) );
  dfnrq1 dff2_bus_ack_reg ( .D(N5433), .CP(n6066), .Q(dff2_bus_ack) );
  dfnrq1 \slave_sel_r_reg[1]  ( .D(N6299), .CP(n6117), .Q(slave_sel_r[1]) );
  dfnrq1 dff_bus_ack_reg ( .D(N5432), .CP(n6066), .Q(dff_bus_ack) );
  dfnrq1 \slave_sel_r_reg[5]  ( .D(N6303), .CP(n6068), .Q(slave_sel_r[5]) );
  dfnrq1 \slave_sel_r_reg[3]  ( .D(N6301), .CP(n6066), .Q(slave_sel_r[3]) );
  dfnrq1 \slave_sel_r_reg[0]  ( .D(N6298), .CP(n6117), .Q(slave_sel_r[0]) );
  dfnrq1 mgmtsoc_vexriscv_transfer_wait_for_ack_reg ( .D(n3401), .CP(n6120), 
        .Q(mgmtsoc_vexriscv_transfer_wait_for_ack) );
  dfnrq1 \slave_sel_r_reg[6]  ( .D(N6304), .CP(n6120), .Q(slave_sel_r[6]) );
  dfnrq1 state_reg ( .D(N6326), .CP(n6117), .Q(state) );
  dfnrq1 mgmtsoc_reset_re_reg ( .D(N5168), .CP(n6120), .Q(mgmtsoc_reset_re) );
  dfnrq1 \spi_master_mosi_storage_reg[0]  ( .D(n4545), .CP(n6120), .Q(
        spi_master_mosi[0]) );
  dfnrq1 \la_out_storage_reg[0]  ( .D(n4480), .CP(n6068), .Q(n134) );
  dfnrq1 \la_out_storage_reg[8]  ( .D(n4472), .CP(n6066), .Q(n126) );
  dfnrq1 \la_out_storage_reg[16]  ( .D(n4464), .CP(n6117), .Q(n118) );
  dfnrq1 \la_out_storage_reg[24]  ( .D(n4456), .CP(n6120), .Q(n110) );
  dfnrq1 \la_out_storage_reg[32]  ( .D(n4448), .CP(n6068), .Q(n102) );
  dfnrq1 \la_out_storage_reg[40]  ( .D(n4440), .CP(n6068), .Q(n94) );
  dfnrq1 \la_out_storage_reg[48]  ( .D(n4432), .CP(n6067), .Q(n86) );
  dfnrq1 \la_out_storage_reg[56]  ( .D(n4424), .CP(n6067), .Q(n78) );
  dfnrq1 \la_out_storage_reg[64]  ( .D(n4416), .CP(n6056), .Q(n70) );
  dfnrq1 \la_out_storage_reg[72]  ( .D(n4408), .CP(n6116), .Q(n62) );
  dfnrq1 \la_out_storage_reg[80]  ( .D(n4400), .CP(n6059), .Q(n54) );
  dfnrq1 \la_out_storage_reg[88]  ( .D(n4392), .CP(n6056), .Q(n46) );
  dfnrq1 \la_out_storage_reg[96]  ( .D(n4384), .CP(n6116), .Q(n38) );
  dfnrq1 \la_out_storage_reg[104]  ( .D(n4376), .CP(n6056), .Q(n30) );
  dfnrq1 \la_out_storage_reg[112]  ( .D(n4368), .CP(n6054), .Q(n22) );
  dfnrq1 \la_out_storage_reg[120]  ( .D(n4360), .CP(n6116), .Q(n14) );
  dfnrq1 \la_oe_storage_reg[0]  ( .D(n4352), .CP(n6059), .Q(csrbank6_oe0_w[0])
         );
  dfnrq1 \la_oe_storage_reg[8]  ( .D(n4344), .CP(n6060), .Q(csrbank6_oe0_w[8])
         );
  dfnrq1 \la_oe_storage_reg[16]  ( .D(n4336), .CP(n6058), .Q(
        csrbank6_oe0_w[16]) );
  dfnrq1 \la_oe_storage_reg[24]  ( .D(n4328), .CP(n6059), .Q(
        csrbank6_oe0_w[24]) );
  dfnrq1 \la_oe_storage_reg[64]  ( .D(n4288), .CP(n6060), .Q(csrbank6_oe2_w[0]) );
  dfnrq1 \la_oe_storage_reg[72]  ( .D(n4280), .CP(n6054), .Q(csrbank6_oe2_w[8]) );
  dfnrq1 \la_oe_storage_reg[80]  ( .D(n4272), .CP(n6054), .Q(
        csrbank6_oe2_w[16]) );
  dfnrq1 \la_oe_storage_reg[88]  ( .D(n4264), .CP(n6054), .Q(
        csrbank6_oe2_w[24]) );
  dfnrq1 \uart_tx_fifo_level0_reg[1]  ( .D(n4040), .CP(n6054), .Q(
        uart_tx_fifo_level0[1]) );
  dfnrq1 \uart_tx_fifo_consume_reg[0]  ( .D(n4052), .CP(n6054), .Q(
        uart_tx_fifo_rdport_adr[0]) );
  dfnrq1 \uart_tx_fifo_consume_reg[1]  ( .D(n4051), .CP(n6054), .Q(
        uart_tx_fifo_rdport_adr[1]) );
  dfnrq1 \uart_tx_fifo_consume_reg[2]  ( .D(n4050), .CP(n6054), .Q(
        uart_tx_fifo_rdport_adr[2]) );
  dfnrq1 \uart_tx_fifo_consume_reg[3]  ( .D(n4049), .CP(n6054), .Q(
        uart_tx_fifo_rdport_adr[3]) );
  dfnrq1 \uart_tx_fifo_level0_reg[0]  ( .D(n4044), .CP(n6062), .Q(
        uart_tx_fifo_level0[0]) );
  dfnrq1 \uart_tx_fifo_level0_reg[4]  ( .D(n4043), .CP(n6054), .Q(
        uart_tx_fifo_level0[4]) );
  dfnrq1 uart_tx_trigger_d_reg ( .D(N5707), .CP(n6060), .Q(uart_tx_trigger_d)
         );
  dfnrq1 \uart_tx_fifo_level0_reg[3]  ( .D(n4042), .CP(n6061), .Q(
        uart_tx_fifo_level0[3]) );
  dfnrq1 \uart_tx_fifo_level0_reg[2]  ( .D(n4041), .CP(n6062), .Q(
        uart_tx_fifo_level0[2]) );
  dfnrq1 uart_tx_fifo_readable_reg ( .D(n3911), .CP(n6054), .Q(
        uart_phy_tx_sink_valid) );
  dfnrq1 rs232phy_rs232phytx_state_reg ( .D(n3904), .CP(n6060), .Q(
        rs232phy_rs232phytx_state) );
  dfnrq1 \uart_phy_tx_phase_reg[5]  ( .D(N3577), .CP(n6061), .Q(
        uart_phy_tx_phase[5]) );
  dfnrq1 \uart_phy_tx_phase_reg[6]  ( .D(N3578), .CP(n6099), .Q(
        uart_phy_tx_phase[6]) );
  dfnrq1 \uart_phy_tx_phase_reg[7]  ( .D(N3579), .CP(n6099), .Q(
        uart_phy_tx_phase[7]) );
  dfnrq1 \uart_phy_tx_phase_reg[8]  ( .D(N3580), .CP(n6028), .Q(
        uart_phy_tx_phase[8]) );
  dfnrq1 \uart_phy_tx_phase_reg[9]  ( .D(N3581), .CP(n6099), .Q(
        uart_phy_tx_phase[9]) );
  dfnrq1 \uart_phy_tx_phase_reg[10]  ( .D(N3582), .CP(n6028), .Q(
        uart_phy_tx_phase[10]) );
  dfnrq1 \uart_phy_tx_phase_reg[11]  ( .D(N3583), .CP(n6028), .Q(
        uart_phy_tx_phase[11]) );
  dfnrq1 \uart_phy_tx_phase_reg[12]  ( .D(N3584), .CP(n6099), .Q(
        uart_phy_tx_phase[12]) );
  dfnrq1 \uart_phy_tx_phase_reg[13]  ( .D(N3585), .CP(n6028), .Q(
        uart_phy_tx_phase[13]) );
  dfnrq1 \uart_phy_tx_phase_reg[14]  ( .D(N3586), .CP(n6055), .Q(
        uart_phy_tx_phase[14]) );
  dfnrq1 \uart_phy_tx_phase_reg[15]  ( .D(N3587), .CP(n6055), .Q(
        uart_phy_tx_phase[15]) );
  dfnrq1 \uart_phy_tx_phase_reg[16]  ( .D(N3588), .CP(n6055), .Q(
        uart_phy_tx_phase[16]) );
  dfnrq1 \uart_phy_tx_phase_reg[17]  ( .D(N3589), .CP(n6055), .Q(
        uart_phy_tx_phase[17]) );
  dfnrq1 \uart_phy_tx_phase_reg[18]  ( .D(N3590), .CP(n6055), .Q(
        uart_phy_tx_phase[18]) );
  dfnrq1 \uart_phy_tx_phase_reg[19]  ( .D(N3591), .CP(n6055), .Q(
        uart_phy_tx_phase[19]) );
  dfnrq1 \uart_phy_tx_phase_reg[20]  ( .D(N3592), .CP(n6055), .Q(
        uart_phy_tx_phase[20]) );
  dfnrq1 \uart_phy_tx_phase_reg[21]  ( .D(N3593), .CP(n6055), .Q(
        uart_phy_tx_phase[21]) );
  dfnrq1 \uart_phy_tx_phase_reg[22]  ( .D(N3594), .CP(n6096), .Q(
        uart_phy_tx_phase[22]) );
  dfnrq1 \uart_phy_tx_phase_reg[23]  ( .D(N3595), .CP(n6124), .Q(
        uart_phy_tx_phase[23]) );
  dfnrq1 \uart_phy_tx_phase_reg[24]  ( .D(N3596), .CP(n6096), .Q(
        uart_phy_tx_phase[24]) );
  dfnrq1 \uart_phy_tx_phase_reg[25]  ( .D(N3597), .CP(n6124), .Q(
        uart_phy_tx_phase[25]) );
  dfnrq1 \uart_phy_tx_phase_reg[26]  ( .D(N3598), .CP(n6096), .Q(
        uart_phy_tx_phase[26]) );
  dfnrq1 \uart_phy_tx_phase_reg[27]  ( .D(N3599), .CP(n6124), .Q(
        uart_phy_tx_phase[27]) );
  dfnrq1 \uart_phy_tx_phase_reg[28]  ( .D(N3600), .CP(n6096), .Q(
        uart_phy_tx_phase[28]) );
  dfnrq1 \uart_phy_tx_phase_reg[29]  ( .D(N3601), .CP(n6124), .Q(
        uart_phy_tx_phase[29]) );
  dfnrq1 \uart_phy_tx_phase_reg[30]  ( .D(N3602), .CP(n6056), .Q(
        uart_phy_tx_phase[30]) );
  dfnrq1 \uart_phy_tx_phase_reg[31]  ( .D(N3603), .CP(n6056), .Q(
        uart_phy_tx_phase[31]) );
  dfnrq1 uart_phy_tx_tick_reg ( .D(N5702), .CP(n6056), .Q(uart_phy_tx_tick) );
  dfnrq1 \uart_phy_tx_count_reg[0]  ( .D(n3903), .CP(n6056), .Q(
        uart_phy_tx_count[0]) );
  dfnrq1 \uart_phy_tx_count_reg[1]  ( .D(n3902), .CP(n6056), .Q(
        uart_phy_tx_count[1]) );
  dfnrq1 \uart_phy_tx_count_reg[2]  ( .D(n3901), .CP(n6056), .Q(
        uart_phy_tx_count[2]) );
  dfnrq1 \uart_phy_tx_count_reg[3]  ( .D(n3900), .CP(n6056), .Q(
        uart_phy_tx_count[3]) );
  dfnrq1 \uart_tx_fifo_produce_reg[0]  ( .D(n4048), .CP(n6128), .Q(
        uart_tx_fifo_produce[0]) );
  dfnrq1 \uart_tx_fifo_produce_reg[1]  ( .D(n4047), .CP(n6025), .Q(
        uart_tx_fifo_produce[1]) );
  dfnrq1 \uart_tx_fifo_produce_reg[2]  ( .D(n4046), .CP(n6128), .Q(
        uart_tx_fifo_produce[2]) );
  dfnrq1 \uart_tx_fifo_produce_reg[3]  ( .D(n4045), .CP(n6025), .Q(
        uart_tx_fifo_produce[3]) );
  dfnrq1 \storage_reg[15][0]  ( .D(n4039), .CP(n6128), .Q(\storage[15][0] ) );
  dfnrq1 \storage_reg[13][0]  ( .D(n4023), .CP(n6025), .Q(\storage[13][0] ) );
  dfnrq1 \storage_reg[11][0]  ( .D(n4007), .CP(n6128), .Q(\storage[11][0] ) );
  dfnrq1 \storage_reg[9][0]  ( .D(n3991), .CP(n6025), .Q(\storage[9][0] ) );
  dfnrq1 \storage_reg[7][0]  ( .D(n3975), .CP(n6057), .Q(\storage[7][0] ) );
  dfnrq1 \storage_reg[5][0]  ( .D(n3959), .CP(n6057), .Q(\storage[5][0] ) );
  dfnrq1 \storage_reg[3][0]  ( .D(n3943), .CP(n6057), .Q(\storage[3][0] ) );
  dfnrq1 \storage_reg[1][0]  ( .D(n3927), .CP(n6057), .Q(\storage[1][0] ) );
  dfnrq1 \storage_reg[14][0]  ( .D(n4031), .CP(n6057), .Q(\storage[14][0] ) );
  dfnrq1 \storage_reg[12][0]  ( .D(n4015), .CP(n6057), .Q(\storage[12][0] ) );
  dfnrq1 \storage_reg[10][0]  ( .D(n3999), .CP(n6057), .Q(\storage[10][0] ) );
  dfnrq1 \storage_reg[8][0]  ( .D(n3983), .CP(n6057), .Q(\storage[8][0] ) );
  dfnrq1 \storage_reg[6][0]  ( .D(n3967), .CP(n6032), .Q(\storage[6][0] ) );
  dfnrq1 \storage_reg[4][0]  ( .D(n3951), .CP(n6022), .Q(\storage[4][0] ) );
  dfnrq1 \storage_reg[2][0]  ( .D(n3935), .CP(n6058), .Q(\storage[2][0] ) );
  dfnrq1 \storage_reg[0][0]  ( .D(n3919), .CP(n6058), .Q(\storage[0][0] ) );
  dfnrq1 \memdat_1_reg[0]  ( .D(n3899), .CP(n6058), .Q(
        uart_tx_fifo_fifo_out_payload_data[0]) );
  dfnrq1 \spimaster_storage_reg[8]  ( .D(n3712), .CP(n6058), .Q(
        spi_master_clk_divider0[8]) );
  dfnrq1 \spi_master_cs_storage_reg[0]  ( .D(n3681), .CP(n6058), .Q(
        csrbank9_cs0_w[0]) );
  dfnrq1 \spi_master_cs_storage_reg[8]  ( .D(n3673), .CP(n6058), .Q(
        csrbank9_cs0_w[8]) );
  dfnrq1 \spi_master_cs_storage_reg[16]  ( .D(n3665), .CP(n6058), .Q(
        csrbank9_cs0_w[16]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[16]  ( .D(N4601), .CP(n6058), .Q(
        interface9_bank_bus_dat_r[16]) );
  dfnrq1 spi_master_control_re_reg ( .D(N5618), .CP(n6058), .Q(
        spi_master_control_re) );
  dfnrq1 \spi_master_control_storage_reg[0]  ( .D(n3664), .CP(n6058), .Q(
        csrbank9_control0_w[0]) );
  dfnrq1 \spimaster_state_reg[0]  ( .D(n3662), .CP(n6046), .Q(
        spimaster_state[0]) );
  dfnrq1 \spimaster_state_reg[1]  ( .D(n3663), .CP(n6046), .Q(
        spimaster_state[1]) );
  dfnrq1 spi_cs_n_reg ( .D(N5589), .CP(n6046), .Q(spi_cs_n) );
  dfnrq1 \spi_master_count_reg[0]  ( .D(n3685), .CP(n6029), .Q(
        spi_master_count[0]) );
  dfnrq1 \spi_master_count_reg[1]  ( .D(n3684), .CP(n6026), .Q(
        spi_master_count[1]) );
  dfnrq1 \spi_master_count_reg[2]  ( .D(n3683), .CP(n6125), .Q(
        spi_master_count[2]) );
  dfnrq1 \spi_master_mosi_sel_reg[0]  ( .D(n3696), .CP(n6046), .Q(
        spi_master_mosi_sel[0]) );
  dfnrq1 \spi_master_mosi_sel_reg[1]  ( .D(n3695), .CP(n6046), .Q(
        spi_master_mosi_sel[1]) );
  dfnrq1 \spi_master_mosi_sel_reg[2]  ( .D(n3694), .CP(n6046), .Q(
        spi_master_mosi_sel[2]) );
  dfnrq1 \spi_master_mosi_data_reg[0]  ( .D(n3693), .CP(n6100), .Q(
        spi_master_mosi_data[0]) );
  dfnrq1 spi_clk_reg ( .D(n3637), .CP(n6023), .Q(spi_clk) );
  dfnrq1 \spi_master_control_storage_reg[8]  ( .D(n3654), .CP(n6058), .Q(
        spi_master_length0[0]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[8]  ( .D(N4593), .CP(n6023), .Q(
        interface9_bank_bus_dat_r[8]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[0]  ( .D(n3559), .CP(n6058), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_len[0]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[8]  ( .D(n3551), .CP(n6023), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_width[0]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[16]  ( .D(n3543), .CP(n6058), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_mask[0]) );
  dfnrq1 mgmtsoc_master_cs_storage_reg ( .D(n3535), .CP(n6023), .Q(
        \litespi_request[1] ) );
  dfnrq1 \mgmtsoc_litespimmap_storage_reg[0]  ( .D(n3534), .CP(n6058), .Q(
        mgmtsoc_litespimmap_spi_dummy_bits[0]) );
  dfnrq1 gpioin5_enable_storage_reg ( .D(n4515), .CP(n6023), .Q(gpioin5_i02)
         );
  dfnrq1 gpioin4_enable_storage_reg ( .D(n4513), .CP(n6059), .Q(gpioin4_i02)
         );
  dfnrq1 gpioin3_enable_storage_reg ( .D(n4511), .CP(n6059), .Q(gpioin3_i02)
         );
  dfnrq1 gpioin2_enable_storage_reg ( .D(n4509), .CP(n6059), .Q(gpioin2_i02)
         );
  dfnrq1 gpioin1_enable_storage_reg ( .D(n4507), .CP(n6059), .Q(gpioin1_i02)
         );
  dfnrq1 gpioin0_enable_storage_reg ( .D(n4505), .CP(n6059), .Q(gpioin0_i02)
         );
  dfnrq1 gpio_out_storage_reg ( .D(n4096), .CP(n6059), .Q(n6130) );
  dfnrq1 \uart_enable_storage_reg[0]  ( .D(n3910), .CP(n6059), .Q(
        csrbank11_ev_enable0_w[0]) );
  dfnrq1 spi_master_loopback_storage_reg ( .D(n3682), .CP(n6059), .Q(
        spi_master_loopback) );
  dfnrq1 mgmtsoc_enable_storage_reg ( .D(n3503), .CP(n6060), .Q(mgmtsoc_zero2)
         );
  dfnrq1 mgmtsoc_pending_re_reg ( .D(N5395), .CP(n6060), .Q(mgmtsoc_pending_re) );
  dfnrq1 mgmtsoc_pending_r_reg ( .D(n3502), .CP(n6060), .Q(mgmtsoc_pending_r)
         );
  dfnrq1 mgmtsoc_update_value_re_reg ( .D(N5358), .CP(n6059), .Q(
        mgmtsoc_update_value_re) );
  dfnrq1 mgmtsoc_update_value_storage_reg ( .D(n3468), .CP(n6043), .Q(
        csrbank10_update_value0_w) );
  dfnrq1 mgmtsoc_en_storage_reg ( .D(n3467), .CP(n6027), .Q(csrbank10_en0_w)
         );
  dfnrq1 \mgmtsoc_reload_storage_reg[0]  ( .D(n3466), .CP(n6127), .Q(
        csrbank10_reload0_w[0]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[8]  ( .D(n3458), .CP(n6127), .Q(
        csrbank10_reload0_w[8]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[16]  ( .D(n3450), .CP(n6031), .Q(
        csrbank10_reload0_w[16]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[24]  ( .D(n3442), .CP(n6030), .Q(
        csrbank10_reload0_w[24]) );
  dfnrq1 \mgmtsoc_load_storage_reg[0]  ( .D(n3434), .CP(n6127), .Q(
        csrbank10_load0_w[0]) );
  dfnrq1 \mgmtsoc_load_storage_reg[8]  ( .D(n3426), .CP(n6030), .Q(
        csrbank10_load0_w[8]) );
  dfnrq1 \mgmtsoc_load_storage_reg[16]  ( .D(n3418), .CP(n6060), .Q(
        csrbank10_load0_w[16]) );
  dfnrq1 \mgmtsoc_load_storage_reg[24]  ( .D(n3410), .CP(n6127), .Q(
        csrbank10_load0_w[24]) );
  dfnrq1 \la_oe_storage_reg[32]  ( .D(n4320), .CP(n6030), .Q(csrbank6_oe1_w[0]) );
  dfnrq1 \la_oe_storage_reg[40]  ( .D(n4312), .CP(n6127), .Q(csrbank6_oe1_w[8]) );
  dfnrq1 \la_oe_storage_reg[48]  ( .D(n4304), .CP(n6030), .Q(
        csrbank6_oe1_w[16]) );
  dfnrq1 \la_oe_storage_reg[56]  ( .D(n4296), .CP(n6061), .Q(
        csrbank6_oe1_w[24]) );
  dfnrq1 \la_ien_storage_reg[0]  ( .D(n4224), .CP(n6127), .Q(
        csrbank6_ien0_w[0]) );
  dfnrq1 \la_ien_storage_reg[8]  ( .D(n4216), .CP(n6031), .Q(
        csrbank6_ien0_w[8]) );
  dfnrq1 \la_ien_storage_reg[16]  ( .D(n4208), .CP(n6127), .Q(
        csrbank6_ien0_w[16]) );
  dfnrq1 \la_ien_storage_reg[24]  ( .D(n4200), .CP(n6127), .Q(
        csrbank6_ien0_w[24]) );
  dfnrq1 gpio_oe_storage_reg ( .D(n4095), .CP(n6062), .Q(csrbank5_oe0_w) );
  dfnrq1 gpioin5_gpioin5_edge_storage_reg ( .D(n4501), .CP(n6030), .Q(
        csrbank18_edge0_w) );
  dfnrq1 gpioin4_gpioin4_edge_storage_reg ( .D(n4498), .CP(n6056), .Q(
        csrbank17_edge0_w) );
  dfnrq1 gpioin3_gpioin3_edge_storage_reg ( .D(n4495), .CP(n6127), .Q(
        csrbank16_edge0_w) );
  dfnrq1 gpioin2_gpioin2_edge_storage_reg ( .D(n4492), .CP(n6031), .Q(
        csrbank15_edge0_w) );
  dfnrq1 gpioin1_gpioin1_edge_storage_reg ( .D(n4489), .CP(n6127), .Q(
        csrbank14_edge0_w) );
  dfnrq1 gpioin0_gpioin0_edge_storage_reg ( .D(n4486), .CP(n6030), .Q(
        csrbank13_edge0_w) );
  dfnrq1 \la_ien_storage_reg[32]  ( .D(n4192), .CP(n6031), .Q(
        csrbank6_ien1_w[0]) );
  dfnrq1 \la_ien_storage_reg[40]  ( .D(n4184), .CP(n6030), .Q(
        csrbank6_ien1_w[8]) );
  dfnrq1 \la_ien_storage_reg[48]  ( .D(n4176), .CP(n6030), .Q(
        csrbank6_ien1_w[16]) );
  dfnrq1 \la_ien_storage_reg[56]  ( .D(n4168), .CP(n6031), .Q(
        csrbank6_ien1_w[24]) );
  dfnrq1 gpio_ien_storage_reg ( .D(n4094), .CP(n6054), .Q(csrbank5_ien0_w) );
  dfnrq1 gpioin5_pending_re_reg ( .D(N6290), .CP(n6031), .Q(gpioin5_pending_re) );
  dfnrq1 gpioin4_pending_re_reg ( .D(N6285), .CP(n6127), .Q(gpioin4_pending_re) );
  dfnrq1 gpioin3_pending_re_reg ( .D(N6280), .CP(n6127), .Q(gpioin3_pending_re) );
  dfnrq1 gpioin2_pending_re_reg ( .D(N6275), .CP(n6031), .Q(gpioin2_pending_re) );
  dfnrq1 gpioin1_pending_re_reg ( .D(N6270), .CP(n6030), .Q(gpioin1_pending_re) );
  dfnrq1 gpioin0_pending_re_reg ( .D(N6265), .CP(n6030), .Q(gpioin0_pending_re) );
  dfnrq1 uart_pending_re_reg ( .D(N5711), .CP(n6030), .Q(uart_pending_re) );
  dfnrq1 gpioin5_pending_r_reg ( .D(n4514), .CP(n6030), .Q(gpioin5_pending_r)
         );
  dfnrq1 gpioin4_pending_r_reg ( .D(n4512), .CP(n6030), .Q(gpioin4_pending_r)
         );
  dfnrq1 gpioin3_pending_r_reg ( .D(n4510), .CP(n6030), .Q(gpioin3_pending_r)
         );
  dfnrq1 gpioin2_pending_r_reg ( .D(n4508), .CP(n6030), .Q(gpioin2_pending_r)
         );
  dfnrq1 gpioin1_pending_r_reg ( .D(n4506), .CP(n6030), .Q(gpioin1_pending_r)
         );
  dfnrq1 gpioin0_pending_r_reg ( .D(n4504), .CP(n6031), .Q(gpioin0_pending_r)
         );
  dfnrq1 \la_oe_storage_reg[96]  ( .D(n4256), .CP(n6031), .Q(csrbank6_oe3_w[0]) );
  dfnrq1 \la_oe_storage_reg[104]  ( .D(n4248), .CP(n6031), .Q(
        csrbank6_oe3_w[8]) );
  dfnrq1 \la_oe_storage_reg[112]  ( .D(n4240), .CP(n6031), .Q(
        csrbank6_oe3_w[16]) );
  dfnrq1 \la_oe_storage_reg[120]  ( .D(n4232), .CP(n6031), .Q(
        csrbank6_oe3_w[24]) );
  dfnrq1 \uart_pending_r_reg[0]  ( .D(n3908), .CP(n6031), .Q(uart_pending_r[0]) );
  dfnrq1 uart_tx_pending_reg ( .D(n3905), .CP(n6031), .Q(
        uart_pending_status[0]) );
  dfnrq1 \user_irq_ena_storage_reg[0]  ( .D(n4484), .CP(n6031), .Q(n6133) );
  dfnrq1 \interface19_bank_bus_dat_r_reg[0]  ( .D(N4995), .CP(n6032), .Q(
        interface19_bank_bus_dat_r[0]) );
  dfnrq1 spi_enabled_storage_reg ( .D(n4481), .CP(n6032), .Q(spi_enabled) );
  dfnrq1 \interface8_bank_bus_dat_r_reg[0]  ( .D(N4516), .CP(n6032), .Q(
        \interface8_bank_bus_dat_r[0] ) );
  dfnrq1 \la_ien_storage_reg[96]  ( .D(n4128), .CP(n6032), .Q(
        csrbank6_ien3_w[0]) );
  dfnrq1 \la_ien_storage_reg[104]  ( .D(n4120), .CP(n6032), .Q(
        csrbank6_ien3_w[8]) );
  dfnrq1 \la_ien_storage_reg[112]  ( .D(n4112), .CP(n6032), .Q(
        csrbank6_ien3_w[16]) );
  dfnrq1 \la_ien_storage_reg[120]  ( .D(n4104), .CP(n6032), .Q(
        csrbank6_ien3_w[24]) );
  dfnrq1 gpio_mode1_storage_reg ( .D(n4092), .CP(n6032), .Q(gpio_mode1_pad) );
  dfnrq1 uart_enabled_storage_reg ( .D(n4091), .CP(n6081), .Q(uart_enabled_o)
         );
  dfnrq1 \interface12_bank_bus_dat_r_reg[0]  ( .D(N4790), .CP(n6036), .Q(
        \interface12_bank_bus_dat_r[0] ) );
  dfnrq1 debug_mode_storage_reg ( .D(n4090), .CP(n6037), .Q(debug_mode) );
  dfnrq1 \interface1_bank_bus_dat_r_reg[0]  ( .D(N4141), .CP(n6048), .Q(
        \interface1_bank_bus_dat_r[0] ) );
  dfnrq1 debug_oeb_storage_reg ( .D(n4089), .CP(n6114), .Q(debug_oeb) );
  dfnrq1 \interface2_bank_bus_dat_r_reg[0]  ( .D(N4152), .CP(n6114), .Q(
        \interface2_bank_bus_dat_r[0] ) );
  dfnrq1 mprj_wb_iena_storage_reg ( .D(n3721), .CP(n6127), .Q(mprj_wb_iena) );
  dfnrq1 \interface7_bank_bus_dat_r_reg[0]  ( .D(N4505), .CP(n6067), .Q(
        \interface7_bank_bus_dat_r[0] ) );
  dfnrq1 \mgmtsoc_litespisdrphycore_storage_reg[0]  ( .D(n3511), .CP(n6067), 
        .Q(mgmtsoc_litespisdrphycore_div[0]) );
  dfnrq1 \interface4_bank_bus_dat_r_reg[0]  ( .D(N4292), .CP(n6126), .Q(
        interface4_bank_bus_dat_r[0]) );
  dfnrq1 gpioin5_gpioin5_mode_storage_reg ( .D(n4500), .CP(n6065), .Q(
        csrbank18_mode0_w) );
  dfnrq1 gpioin5_gpioin5_trigger_d_reg ( .D(N6247), .CP(n6035), .Q(
        gpioin5_gpioin5_trigger_d) );
  dfnrq1 gpioin5_gpioin5_pending_reg ( .D(n4502), .CP(n6118), .Q(gpioin5_i01)
         );
  dfnrq1 \interface18_bank_bus_dat_r_reg[0]  ( .D(N4982), .CP(n6063), .Q(
        \interface18_bank_bus_dat_r[0] ) );
  dfnrq1 gpioin4_gpioin4_mode_storage_reg ( .D(n4497), .CP(n6126), .Q(
        csrbank17_mode0_w) );
  dfnrq1 gpioin4_gpioin4_trigger_d_reg ( .D(N6239), .CP(n6034), .Q(
        gpioin4_gpioin4_trigger_d) );
  dfnrq1 gpioin4_gpioin4_pending_reg ( .D(n4499), .CP(n6125), .Q(gpioin4_i01)
         );
  dfnrq1 \interface17_bank_bus_dat_r_reg[0]  ( .D(N4950), .CP(n6025), .Q(
        \interface17_bank_bus_dat_r[0] ) );
  dfnrq1 gpioin3_gpioin3_mode_storage_reg ( .D(n4494), .CP(n6126), .Q(
        csrbank16_mode0_w) );
  dfnrq1 gpioin3_gpioin3_trigger_d_reg ( .D(N6231), .CP(n6024), .Q(
        gpioin3_gpioin3_trigger_d) );
  dfnrq1 gpioin3_gpioin3_pending_reg ( .D(n4496), .CP(n6126), .Q(gpioin3_i01)
         );
  dfnrq1 \interface16_bank_bus_dat_r_reg[0]  ( .D(N4918), .CP(n6067), .Q(
        \interface16_bank_bus_dat_r[0] ) );
  dfnrq1 gpioin2_gpioin2_mode_storage_reg ( .D(n4491), .CP(n6035), .Q(
        csrbank15_mode0_w) );
  dfnrq1 gpioin2_gpioin2_trigger_d_reg ( .D(N6223), .CP(n6050), .Q(
        gpioin2_gpioin2_trigger_d) );
  dfnrq1 gpioin2_gpioin2_pending_reg ( .D(n4493), .CP(n6047), .Q(gpioin2_i01)
         );
  dfnrq1 \interface15_bank_bus_dat_r_reg[0]  ( .D(N4886), .CP(n6034), .Q(
        \interface15_bank_bus_dat_r[0] ) );
  dfnrq1 gpioin1_gpioin1_mode_storage_reg ( .D(n4488), .CP(n6126), .Q(
        csrbank14_mode0_w) );
  dfnrq1 gpioin1_gpioin1_trigger_d_reg ( .D(N6215), .CP(n6114), .Q(
        gpioin1_gpioin1_trigger_d) );
  dfnrq1 gpioin1_gpioin1_pending_reg ( .D(n4490), .CP(n6035), .Q(gpioin1_i01)
         );
  dfnrq1 \interface14_bank_bus_dat_r_reg[0]  ( .D(N4854), .CP(n6034), .Q(
        \interface14_bank_bus_dat_r[0] ) );
  dfnrq1 gpioin0_gpioin0_mode_storage_reg ( .D(n4485), .CP(n6100), .Q(
        csrbank13_mode0_w) );
  dfnrq1 gpioin0_gpioin0_trigger_d_reg ( .D(N6207), .CP(n6033), .Q(
        gpioin0_gpioin0_trigger_d) );
  dfnrq1 gpioin0_gpioin0_pending_reg ( .D(n4487), .CP(n6056), .Q(gpioin0_i01)
         );
  dfnrq1 \interface13_bank_bus_dat_r_reg[0]  ( .D(N4822), .CP(n6126), .Q(
        \interface13_bank_bus_dat_r[0] ) );
  dfnrq1 \la_ien_storage_reg[64]  ( .D(n4160), .CP(n6126), .Q(
        csrbank6_ien2_w[0]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[0]  ( .D(N4463), .CP(n6116), .Q(
        interface6_bank_bus_dat_r[0]) );
  dfnrq1 \la_ien_storage_reg[72]  ( .D(n4152), .CP(n6034), .Q(
        csrbank6_ien2_w[8]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[8]  ( .D(N4471), .CP(n6126), .Q(
        interface6_bank_bus_dat_r[8]) );
  dfnrq1 \la_ien_storage_reg[80]  ( .D(n4144), .CP(n6035), .Q(
        csrbank6_ien2_w[16]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[16]  ( .D(N4479), .CP(n6033), .Q(
        interface6_bank_bus_dat_r[16]) );
  dfnrq1 \la_ien_storage_reg[88]  ( .D(n4136), .CP(n6033), .Q(
        csrbank6_ien2_w[24]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[24]  ( .D(N4487), .CP(n6033), .Q(
        interface6_bank_bus_dat_r[24]) );
  dfnrq1 gpio_mode0_storage_reg ( .D(n4093), .CP(n6033), .Q(gpio_mode0_pad) );
  dfnrq1 \interface5_bank_bus_dat_r_reg[0]  ( .D(N4331), .CP(n6033), .Q(
        \interface5_bank_bus_dat_r[0] ) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[0]  ( .D(n3327), .CP(n6033), .Q(
        csrbank0_scratch0_w[0]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[8]  ( .D(n3319), .CP(n6033), .Q(
        csrbank0_scratch0_w[8]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[8]  ( .D(N4107), .CP(n6033), .Q(
        interface0_bank_bus_dat_r[8]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[16]  ( .D(n3311), .CP(n6071), .Q(
        csrbank0_scratch0_w[16]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[16]  ( .D(N4115), .CP(n6034), .Q(
        interface0_bank_bus_dat_r[16]) );
  dfnrq1 \mgmtsoc_reset_storage_reg[0]  ( .D(n3295), .CP(n6065), .Q(
        csrbank0_reset0_w[0]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[0]  ( .D(N4099), .CP(n6064), .Q(
        interface0_bank_bus_dat_r[0]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[29]  ( .D(n3192), .CP(n6126), .Q(
        mgmtsoc_litespimmap_burst_adr[29]) );
  dfnrq1 litespi_grant_reg ( .D(n4503), .CP(n6027), .Q(litespi_tx_mux_sel) );
  dfnrq1 \mgmtsoc_litespisdrphycore_count_reg[1]  ( .D(n3513), .CP(n6034), .Q(
        mgmtsoc_litespisdrphycore_count[1]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_count_reg[3]  ( .D(n3515), .CP(n6028), .Q(
        mgmtsoc_litespisdrphycore_count[3]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_count_reg[0]  ( .D(n3516), .CP(n6096), .Q(
        mgmtsoc_litespisdrphycore_count[0]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_count_reg[2]  ( .D(n3514), .CP(n6025), .Q(
        mgmtsoc_litespisdrphycore_count[2]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_cnt_reg[7]  ( .D(n3120), .CP(n6057), 
        .Q(mgmtsoc_litespisdrphycore_sr_cnt[7]) );
  dfnrq1 \litespiphy_state_reg[1]  ( .D(N6249), .CP(n6056), .Q(
        litespiphy_state[1]) );
  dfnrq1 \litespi_state_reg[1]  ( .D(N6253), .CP(n6023), .Q(litespi_state[1])
         );
  dfnrq1 \dbg_uart_data_reg[31]  ( .D(n3252), .CP(n6026), .Q(
        dbg_uart_wishbone_dat_w[31]) );
  dfnrq1 \la_out_storage_reg[31]  ( .D(n4449), .CP(n6112), .Q(n103) );
  dfnrq1 \la_out_storage_reg[63]  ( .D(n4417), .CP(n6128), .Q(n71) );
  dfnrq1 \la_out_storage_reg[95]  ( .D(n4385), .CP(n6112), .Q(n39) );
  dfnrq1 \la_out_storage_reg[127]  ( .D(n4353), .CP(n6032), .Q(n7) );
  dfnrq1 \la_oe_storage_reg[31]  ( .D(n4321), .CP(n6112), .Q(
        csrbank6_oe0_w[31]) );
  dfnrq1 \la_oe_storage_reg[63]  ( .D(n4289), .CP(n6096), .Q(
        csrbank6_oe1_w[31]) );
  dfnrq1 \la_oe_storage_reg[95]  ( .D(n4257), .CP(n6112), .Q(
        csrbank6_oe2_w[31]) );
  dfnrq1 \la_oe_storage_reg[127]  ( .D(n4225), .CP(n6089), .Q(
        csrbank6_oe3_w[31]) );
  dfnrq1 \la_ien_storage_reg[31]  ( .D(n4193), .CP(n6112), .Q(
        csrbank6_ien0_w[31]) );
  dfnrq1 \la_ien_storage_reg[63]  ( .D(n4161), .CP(n6088), .Q(
        csrbank6_ien1_w[31]) );
  dfnrq1 \la_ien_storage_reg[95]  ( .D(n4129), .CP(n6112), .Q(
        csrbank6_ien2_w[31]) );
  dfnrq1 \la_ien_storage_reg[127]  ( .D(n4097), .CP(n6101), .Q(
        csrbank6_ien3_w[31]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[31]  ( .D(N4494), .CP(n6112), .Q(
        interface6_bank_bus_dat_r[31]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[31]  ( .D(n3435), .CP(n6101), .Q(
        csrbank10_reload0_w[31]) );
  dfnrq1 \mgmtsoc_load_storage_reg[31]  ( .D(n3403), .CP(n6112), .Q(
        csrbank10_load0_w[31]) );
  dfnrq1 \mgmtsoc_value_reg[31]  ( .D(N5431), .CP(n6044), .Q(mgmtsoc_value[31]) );
  dfnrq1 mgmtsoc_zero_trigger_d_reg ( .D(N5394), .CP(n6112), .Q(
        mgmtsoc_zero_trigger_d) );
  dfnrq1 \mgmtsoc_value_reg[0]  ( .D(N5400), .CP(n6029), .Q(mgmtsoc_value[0])
         );
  dfnrq1 \mgmtsoc_value_status_reg[0]  ( .D(n3500), .CP(n6112), .Q(
        csrbank10_value_w[0]) );
  dfnrq1 \mgmtsoc_value_reg[8]  ( .D(N5408), .CP(n6097), .Q(mgmtsoc_value[8])
         );
  dfnrq1 \mgmtsoc_value_status_reg[8]  ( .D(n3492), .CP(n6112), .Q(
        csrbank10_value_w[8]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[8]  ( .D(N4702), .CP(n6098), .Q(
        interface10_bank_bus_dat_r[8]) );
  dfnrq1 \mgmtsoc_value_reg[16]  ( .D(N5416), .CP(n6112), .Q(mgmtsoc_value[16]) );
  dfnrq1 \mgmtsoc_value_status_reg[16]  ( .D(n3484), .CP(n6074), .Q(
        csrbank10_value_w[16]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[16]  ( .D(N4710), .CP(n6022), .Q(
        interface10_bank_bus_dat_r[16]) );
  dfnrq1 \mgmtsoc_value_reg[24]  ( .D(N5424), .CP(n6022), .Q(mgmtsoc_value[24]) );
  dfnrq1 \mgmtsoc_value_status_reg[24]  ( .D(n3476), .CP(n6022), .Q(
        csrbank10_value_w[24]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[24]  ( .D(N4718), .CP(n6022), .Q(
        interface10_bank_bus_dat_r[24]) );
  dfnrq1 \mgmtsoc_value_reg[30]  ( .D(N5430), .CP(n6022), .Q(mgmtsoc_value[30]) );
  dfnrq1 \mgmtsoc_value_status_reg[30]  ( .D(n3470), .CP(n6022), .Q(
        csrbank10_value_w[30]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[30]  ( .D(N4724), .CP(n6022), .Q(
        interface10_bank_bus_dat_r[30]) );
  dfnrq1 \dbg_uart_data_reg[30]  ( .D(n3253), .CP(n6022), .Q(
        dbg_uart_wishbone_dat_w[30]) );
  dfnrq1 \dbg_uart_data_reg[29]  ( .D(n3254), .CP(n6023), .Q(
        dbg_uart_wishbone_dat_w[29]) );
  dfnrq1 \dbg_uart_data_reg[28]  ( .D(n3255), .CP(n6023), .Q(
        dbg_uart_wishbone_dat_w[28]) );
  dfnrq1 \dbg_uart_data_reg[11]  ( .D(n3272), .CP(n6023), .Q(
        dbg_uart_wishbone_dat_w[11]) );
  dfnrq1 \la_out_storage_reg[11]  ( .D(n4469), .CP(n6023), .Q(n123) );
  dfnrq1 \la_out_storage_reg[43]  ( .D(n4437), .CP(n6023), .Q(n91) );
  dfnrq1 \la_out_storage_reg[75]  ( .D(n4405), .CP(n6023), .Q(n59) );
  dfnrq1 \la_out_storage_reg[107]  ( .D(n4373), .CP(n6023), .Q(n27) );
  dfnrq1 \la_oe_storage_reg[11]  ( .D(n4341), .CP(n6023), .Q(
        csrbank6_oe0_w[11]) );
  dfnrq1 \la_oe_storage_reg[43]  ( .D(n4309), .CP(n6024), .Q(
        csrbank6_oe1_w[11]) );
  dfnrq1 \la_oe_storage_reg[75]  ( .D(n4277), .CP(n6024), .Q(
        csrbank6_oe2_w[11]) );
  dfnrq1 \la_oe_storage_reg[107]  ( .D(n4245), .CP(n6024), .Q(
        csrbank6_oe3_w[11]) );
  dfnrq1 \la_ien_storage_reg[11]  ( .D(n4213), .CP(n6024), .Q(
        csrbank6_ien0_w[11]) );
  dfnrq1 \la_ien_storage_reg[43]  ( .D(n4181), .CP(n6024), .Q(
        csrbank6_ien1_w[11]) );
  dfnrq1 \la_ien_storage_reg[75]  ( .D(n4149), .CP(n6024), .Q(
        csrbank6_ien2_w[11]) );
  dfnrq1 \la_ien_storage_reg[107]  ( .D(n4117), .CP(n6024), .Q(
        csrbank6_ien3_w[11]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[11]  ( .D(N4474), .CP(n6024), .Q(
        interface6_bank_bus_dat_r[11]) );
  dfnrq1 \spimaster_storage_reg[11]  ( .D(n3709), .CP(n6025), .Q(
        spi_master_clk_divider0[11]) );
  dfnrq1 \spi_master_cs_storage_reg[11]  ( .D(n3670), .CP(n6025), .Q(
        csrbank9_cs0_w[11]) );
  dfnrq1 \spi_master_control_storage_reg[11]  ( .D(n3651), .CP(n6025), .Q(
        spi_master_length0[3]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[11]  ( .D(N4596), .CP(n6025), .Q(
        interface9_bank_bus_dat_r[11]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[11]  ( .D(n3548), .CP(n6025), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_width[3]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_width_reg[3]  ( .D(n3561), 
        .CP(n6025), .Q(mgmtsoc_port_master_user_port_sink_payload_width[3]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[31]  ( .D(n3160), .CP(n6025), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[31]) );
  dfnrq1 \dbg_uart_data_reg[7]  ( .D(n3276), .CP(n6025), .Q(
        dbg_uart_wishbone_dat_w[7]) );
  dfnrq1 \spi_master_mosi_storage_reg[7]  ( .D(n4538), .CP(n6026), .Q(
        spi_master_mosi[7]) );
  dfnrq1 \spi_master_mosi_data_reg[7]  ( .D(n3686), .CP(n6026), .Q(
        spi_master_mosi_data[7]) );
  dfnrq1 \la_out_storage_reg[7]  ( .D(n4473), .CP(n6026), .Q(n127) );
  dfnrq1 \la_out_storage_reg[39]  ( .D(n4441), .CP(n6026), .Q(n95) );
  dfnrq1 \la_out_storage_reg[71]  ( .D(n4409), .CP(n6026), .Q(n63) );
  dfnrq1 \la_out_storage_reg[103]  ( .D(n4377), .CP(n6026), .Q(n31) );
  dfnrq1 \la_oe_storage_reg[7]  ( .D(n4345), .CP(n6026), .Q(csrbank6_oe0_w[7])
         );
  dfnrq1 \la_oe_storage_reg[39]  ( .D(n4313), .CP(n6027), .Q(csrbank6_oe1_w[7]) );
  dfnrq1 \la_oe_storage_reg[71]  ( .D(n4281), .CP(n6027), .Q(csrbank6_oe2_w[7]) );
  dfnrq1 \la_oe_storage_reg[103]  ( .D(n4249), .CP(n6027), .Q(
        csrbank6_oe3_w[7]) );
  dfnrq1 \la_ien_storage_reg[7]  ( .D(n4217), .CP(n6027), .Q(
        csrbank6_ien0_w[7]) );
  dfnrq1 \la_ien_storage_reg[39]  ( .D(n4185), .CP(n6027), .Q(
        csrbank6_ien1_w[7]) );
  dfnrq1 \la_ien_storage_reg[71]  ( .D(n4153), .CP(n6027), .Q(
        csrbank6_ien2_w[7]) );
  dfnrq1 \la_ien_storage_reg[103]  ( .D(n4121), .CP(n6027), .Q(
        csrbank6_ien3_w[7]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[7]  ( .D(N4470), .CP(n6027), .Q(
        interface6_bank_bus_dat_r[7]) );
  dfnrq1 \storage_reg[15][7]  ( .D(n4032), .CP(n6028), .Q(\storage[15][7] ) );
  dfnrq1 \storage_reg[14][7]  ( .D(n4024), .CP(n6028), .Q(\storage[14][7] ) );
  dfnrq1 \storage_reg[13][7]  ( .D(n4016), .CP(n6028), .Q(\storage[13][7] ) );
  dfnrq1 \storage_reg[12][7]  ( .D(n4008), .CP(n6028), .Q(\storage[12][7] ) );
  dfnrq1 \storage_reg[11][7]  ( .D(n4000), .CP(n6028), .Q(\storage[11][7] ) );
  dfnrq1 \storage_reg[10][7]  ( .D(n3992), .CP(n6028), .Q(\storage[10][7] ) );
  dfnrq1 \storage_reg[9][7]  ( .D(n3984), .CP(n6028), .Q(\storage[9][7] ) );
  dfnrq1 \storage_reg[8][7]  ( .D(n3976), .CP(n6028), .Q(\storage[8][7] ) );
  dfnrq1 \storage_reg[7][7]  ( .D(n3968), .CP(n6029), .Q(\storage[7][7] ) );
  dfnrq1 \storage_reg[6][7]  ( .D(n3960), .CP(n6029), .Q(\storage[6][7] ) );
  dfnrq1 \storage_reg[5][7]  ( .D(n3952), .CP(n6029), .Q(\storage[5][7] ) );
  dfnrq1 \storage_reg[4][7]  ( .D(n3944), .CP(n6029), .Q(\storage[4][7] ) );
  dfnrq1 \storage_reg[3][7]  ( .D(n3936), .CP(n6029), .Q(\storage[3][7] ) );
  dfnrq1 \storage_reg[2][7]  ( .D(n3928), .CP(n6029), .Q(\storage[2][7] ) );
  dfnrq1 \storage_reg[1][7]  ( .D(n3920), .CP(n6029), .Q(\storage[1][7] ) );
  dfnrq1 \storage_reg[0][7]  ( .D(n3912), .CP(n6029), .Q(\storage[0][7] ) );
  dfnrq1 \memdat_1_reg[7]  ( .D(n3898), .CP(n6036), .Q(
        uart_tx_fifo_fifo_out_payload_data[7]) );
  dfnrq1 \uart_phy_tx_data_reg[7]  ( .D(n3884), .CP(n6044), .Q(
        uart_phy_tx_data[7]) );
  dfnrq1 \spimaster_storage_reg[7]  ( .D(n3713), .CP(n6045), .Q(
        spi_master_clk_divider0[7]) );
  dfnrq1 \spi_master_cs_storage_reg[7]  ( .D(n3674), .CP(n6112), .Q(
        csrbank9_cs0_w[7]) );
  dfnrq1 \spi_master_control_storage_reg[7]  ( .D(n3655), .CP(n6029), .Q(
        csrbank9_control0_w[7]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[7]  ( .D(n3552), .CP(n6051), 
        .Q(mgmtsoc_master_len[7]) );
  dfnrq1 \mgmtsoc_litespimmap_storage_reg[7]  ( .D(n3527), .CP(n6055), .Q(
        mgmtsoc_litespimmap_spi_dummy_bits[7]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_storage_reg[7]  ( .D(n3504), .CP(n6075), 
        .Q(mgmtsoc_litespisdrphycore_div[7]) );
  dfnrq1 \interface4_bank_bus_dat_r_reg[7]  ( .D(N4299), .CP(n6050), .Q(
        interface4_bank_bus_dat_r[7]) );
  dfnrq1 mgmtsoc_litespisdrphycore_posedge_reg_reg ( .D(N5453), .CP(n6050), 
        .Q(mgmtsoc_litespisdrphycore_posedge_reg) );
  dfnrq1 mgmtsoc_litespisdrphycore_posedge_reg2_reg ( .D(N5454), .CP(n6052), 
        .Q(mgmtsoc_litespisdrphycore_posedge_reg2) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[0]  ( .D(n3190), .CP(n6051), .Q(
        mgmtsoc_litespisdrphycore_source_payload_data[0]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[29]  ( .D(n3161), .CP(n6055), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[29]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[30]  ( .D(n3191), .CP(n6053), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[30]) );
  dfnrq1 \dbg_uart_data_reg[6]  ( .D(n3277), .CP(n6053), .Q(
        dbg_uart_wishbone_dat_w[6]) );
  dfnrq1 \spi_master_mosi_storage_reg[6]  ( .D(n4539), .CP(n6127), .Q(
        spi_master_mosi[6]) );
  dfnrq1 \spi_master_mosi_data_reg[6]  ( .D(n3687), .CP(n6030), .Q(
        spi_master_mosi_data[6]) );
  dfnrq1 \la_out_storage_reg[6]  ( .D(n4474), .CP(n6028), .Q(n128) );
  dfnrq1 \la_out_storage_reg[38]  ( .D(n4442), .CP(n6031), .Q(n96) );
  dfnrq1 \la_out_storage_reg[70]  ( .D(n4410), .CP(n6127), .Q(n64) );
  dfnrq1 \la_out_storage_reg[102]  ( .D(n4378), .CP(n6031), .Q(n32) );
  dfnrq1 \la_oe_storage_reg[6]  ( .D(n4346), .CP(n6127), .Q(csrbank6_oe0_w[6])
         );
  dfnrq1 \la_oe_storage_reg[38]  ( .D(n4314), .CP(n6115), .Q(csrbank6_oe1_w[6]) );
  dfnrq1 \la_oe_storage_reg[70]  ( .D(n4282), .CP(n6115), .Q(csrbank6_oe2_w[6]) );
  dfnrq1 \la_oe_storage_reg[102]  ( .D(n4250), .CP(n6030), .Q(
        csrbank6_oe3_w[6]) );
  dfnrq1 \la_ien_storage_reg[6]  ( .D(n4218), .CP(n6062), .Q(
        csrbank6_ien0_w[6]) );
  dfnrq1 \la_ien_storage_reg[38]  ( .D(n4186), .CP(n6127), .Q(
        csrbank6_ien1_w[6]) );
  dfnrq1 \la_ien_storage_reg[70]  ( .D(n4154), .CP(n6127), .Q(
        csrbank6_ien2_w[6]) );
  dfnrq1 \la_ien_storage_reg[102]  ( .D(n4122), .CP(n6030), .Q(
        csrbank6_ien3_w[6]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[6]  ( .D(N4469), .CP(n6127), .Q(
        interface6_bank_bus_dat_r[6]) );
  dfnrq1 \storage_reg[15][6]  ( .D(n4033), .CP(n6031), .Q(\storage[15][6] ) );
  dfnrq1 \storage_reg[14][6]  ( .D(n4025), .CP(n6041), .Q(\storage[14][6] ) );
  dfnrq1 \storage_reg[13][6]  ( .D(n4017), .CP(n6049), .Q(\storage[13][6] ) );
  dfnrq1 \storage_reg[12][6]  ( .D(n4009), .CP(n6087), .Q(\storage[12][6] ) );
  dfnrq1 \storage_reg[11][6]  ( .D(n4001), .CP(n6113), .Q(\storage[11][6] ) );
  dfnrq1 \storage_reg[10][6]  ( .D(n3993), .CP(n6040), .Q(\storage[10][6] ) );
  dfnrq1 \storage_reg[9][6]  ( .D(n3985), .CP(n6087), .Q(\storage[9][6] ) );
  dfnrq1 \storage_reg[8][6]  ( .D(n3977), .CP(n6113), .Q(\storage[8][6] ) );
  dfnrq1 \storage_reg[7][6]  ( .D(n3969), .CP(n6042), .Q(\storage[7][6] ) );
  dfnrq1 \storage_reg[6][6]  ( .D(n3961), .CP(n6049), .Q(\storage[6][6] ) );
  dfnrq1 \storage_reg[5][6]  ( .D(n3953), .CP(n6042), .Q(\storage[5][6] ) );
  dfnrq1 \storage_reg[4][6]  ( .D(n3945), .CP(n6043), .Q(\storage[4][6] ) );
  dfnrq1 \storage_reg[3][6]  ( .D(n3937), .CP(n6049), .Q(\storage[3][6] ) );
  dfnrq1 \storage_reg[2][6]  ( .D(n3929), .CP(n6113), .Q(\storage[2][6] ) );
  dfnrq1 \storage_reg[1][6]  ( .D(n3921), .CP(n6042), .Q(\storage[1][6] ) );
  dfnrq1 \storage_reg[0][6]  ( .D(n3913), .CP(n6042), .Q(\storage[0][6] ) );
  dfnrq1 \memdat_1_reg[6]  ( .D(n3897), .CP(n6043), .Q(
        uart_tx_fifo_fifo_out_payload_data[6]) );
  dfnrq1 \uart_phy_tx_data_reg[6]  ( .D(n3885), .CP(n6049), .Q(
        uart_phy_tx_data[6]) );
  dfnrq1 \spimaster_storage_reg[6]  ( .D(n3714), .CP(n6040), .Q(
        spi_master_clk_divider0[6]) );
  dfnrq1 \spi_master_cs_storage_reg[6]  ( .D(n3675), .CP(n6087), .Q(
        csrbank9_cs0_w[6]) );
  dfnrq1 \spi_master_control_storage_reg[6]  ( .D(n3656), .CP(n6113), .Q(
        csrbank9_control0_w[6]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[6]  ( .D(n3553), .CP(n6040), 
        .Q(mgmtsoc_master_len[6]) );
  dfnrq1 \mgmtsoc_litespimmap_storage_reg[6]  ( .D(n3528), .CP(n6087), .Q(
        mgmtsoc_litespimmap_spi_dummy_bits[6]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_storage_reg[6]  ( .D(n3505), .CP(n6113), 
        .Q(mgmtsoc_litespisdrphycore_div[6]) );
  dfnrq1 \interface4_bank_bus_dat_r_reg[6]  ( .D(N4298), .CP(n6042), .Q(
        interface4_bank_bus_dat_r[6]) );
  dfnrq1 \litespi_state_reg[3]  ( .D(N6255), .CP(n6043), .Q(litespi_state[3])
         );
  dfnrq1 \litespi_state_reg[2]  ( .D(N6254), .CP(n6049), .Q(litespi_state[2])
         );
  dfnrq1 \litespi_state_reg[0]  ( .D(N6252), .CP(n6040), .Q(litespi_state[0])
         );
  dfnrq1 \litespiphy_state_reg[0]  ( .D(N6248), .CP(n6087), .Q(
        litespiphy_state[0]) );
  dfnrq1 mgmtsoc_master_rx_fifo_source_valid_reg ( .D(n3636), .CP(n6125), .Q(
        \mgmtsoc_master_status_status[1] ) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[0]  ( .D(n3635), .CP(
        n6046), .Q(mgmtsoc_master_rxtx_w[0]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[29]  ( .D(n3606), 
        .CP(n6112), .Q(mgmtsoc_master_rxtx_w[29]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[29]  ( .D(N4272), .CP(n6046), .Q(
        interface3_bank_bus_dat_r[29]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[30]  ( .D(n3605), 
        .CP(n6089), .Q(mgmtsoc_master_rxtx_w[30]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[30]  ( .D(N4273), .CP(n6046), .Q(
        interface3_bank_bus_dat_r[30]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[31]  ( .D(n3604), 
        .CP(n6094), .Q(mgmtsoc_master_rxtx_w[31]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[31]  ( .D(N4274), .CP(n6046), .Q(
        interface3_bank_bus_dat_r[31]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_cnt_reg[0]  ( .D(N5443), .CP(n6114), .Q(
        mgmtsoc_litespisdrphycore_cnt[0]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_cnt_reg[1]  ( .D(N5444), .CP(n6037), .Q(
        mgmtsoc_litespisdrphycore_cnt[1]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_cnt_reg[2]  ( .D(N5445), .CP(n6114), .Q(
        mgmtsoc_litespisdrphycore_cnt[2]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_cnt_reg[3]  ( .D(N5446), .CP(n6038), .Q(
        mgmtsoc_litespisdrphycore_cnt[3]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_cnt_reg[4]  ( .D(N5447), .CP(n6048), .Q(
        mgmtsoc_litespisdrphycore_cnt[4]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_cnt_reg[5]  ( .D(N5448), .CP(n6036), .Q(
        mgmtsoc_litespisdrphycore_cnt[5]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_cnt_reg[6]  ( .D(N5449), .CP(n6037), .Q(
        mgmtsoc_litespisdrphycore_cnt[6]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_cnt_reg[7]  ( .D(N5450), .CP(n6038), .Q(
        mgmtsoc_litespisdrphycore_cnt[7]) );
  dfnrq1 mgmtsoc_litespisdrphycore_clk_reg ( .D(n3512), .CP(n6040), .Q(
        mgmtsoc_litespisdrphycore_clk) );
  dfnrq1 \mgmtsoc_litespimmap_count_reg[0]  ( .D(n3526), .CP(n6043), .Q(
        mgmtsoc_litespimmap_count[0]) );
  dfnrq1 \mgmtsoc_litespimmap_count_reg[7]  ( .D(n3524), .CP(n6049), .Q(
        mgmtsoc_litespimmap_count[7]) );
  dfnrq1 \mgmtsoc_litespimmap_count_reg[6]  ( .D(n3523), .CP(n6113), .Q(
        mgmtsoc_litespimmap_count[6]) );
  dfnrq1 \mgmtsoc_litespimmap_count_reg[5]  ( .D(n3522), .CP(n6042), .Q(
        mgmtsoc_litespimmap_count[5]) );
  dfnrq1 \mgmtsoc_litespimmap_count_reg[4]  ( .D(n3521), .CP(n6090), .Q(
        mgmtsoc_litespimmap_count[4]) );
  dfnrq1 \mgmtsoc_litespimmap_count_reg[3]  ( .D(n3520), .CP(n6091), .Q(
        mgmtsoc_litespimmap_count[3]) );
  dfnrq1 \mgmtsoc_litespimmap_count_reg[2]  ( .D(n3519), .CP(n6093), .Q(
        mgmtsoc_litespimmap_count[2]) );
  dfnrq1 \mgmtsoc_litespimmap_count_reg[1]  ( .D(n3518), .CP(n6040), .Q(
        mgmtsoc_litespimmap_count[1]) );
  dfnrq1 \mgmtsoc_litespimmap_count_reg[8]  ( .D(n3525), .CP(n6040), .Q(
        mgmtsoc_litespimmap_count[8]) );
  dfnrq1 mgmtsoc_litespimmap_burst_cs_reg ( .D(n3517), .CP(n6040), .Q(
        mgmtsoc_litespimmap_burst_cs) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[0]  ( .D(N4243), .CP(n6040), .Q(
        interface3_bank_bus_dat_r[0]) );
  dfnrq1 mgmtsoc_master_tx_fifo_source_valid_reg ( .D(n3603), .CP(n6040), .Q(
        mgmtsoc_port_master_user_port_sink_valid) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[0]  ( .D(n3602), .CP(
        n6040), .Q(mgmtsoc_port_master_user_port_sink_payload_data[0]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[6]  ( .D(n3596), .CP(
        n6040), .Q(mgmtsoc_port_master_user_port_sink_payload_data[6]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[7]  ( .D(n3595), .CP(
        n6040), .Q(mgmtsoc_port_master_user_port_sink_payload_data[7]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[8]  ( .D(n3594), .CP(
        n6041), .Q(mgmtsoc_port_master_user_port_sink_payload_data[8]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[11]  ( .D(n3591), 
        .CP(n6041), .Q(mgmtsoc_port_master_user_port_sink_payload_data[11]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[16]  ( .D(n3586), 
        .CP(n6041), .Q(mgmtsoc_port_master_user_port_sink_payload_data[16]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[24]  ( .D(n3578), 
        .CP(n6041), .Q(mgmtsoc_port_master_user_port_sink_payload_data[24]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[31]  ( .D(n3571), 
        .CP(n6041), .Q(mgmtsoc_port_master_user_port_sink_payload_data[31]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_len_reg[0]  ( .D(n3570), .CP(
        n6041), .Q(mgmtsoc_port_master_user_port_sink_payload_len[0]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_width_reg[0]  ( .D(n3564), 
        .CP(n6041), .Q(mgmtsoc_port_master_user_port_sink_payload_width[0]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_width_reg[2]  ( .D(n3562), 
        .CP(n6042), .Q(mgmtsoc_port_master_user_port_sink_payload_width[2]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[1]  ( .D(n3189), .CP(n6042), .Q(
        mgmtsoc_litespisdrphycore_source_payload_data[1]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[1]  ( .D(n3634), .CP(
        n6042), .Q(mgmtsoc_master_rxtx_w[1]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[2]  ( .D(n3188), .CP(n6042), .Q(
        mgmtsoc_litespisdrphycore_source_payload_data[2]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[2]  ( .D(n3633), .CP(
        n6042), .Q(mgmtsoc_master_rxtx_w[2]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[3]  ( .D(n3187), .CP(n6042), .Q(
        mgmtsoc_litespisdrphycore_source_payload_data[3]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[3]  ( .D(n3632), .CP(
        n6042), .Q(mgmtsoc_master_rxtx_w[3]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[4]  ( .D(n3186), .CP(n6042), .Q(
        mgmtsoc_litespisdrphycore_source_payload_data[4]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[4]  ( .D(n3631), .CP(
        n6091), .Q(mgmtsoc_master_rxtx_w[4]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[5]  ( .D(n3185), .CP(n6125), .Q(
        mgmtsoc_litespisdrphycore_source_payload_data[5]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[5]  ( .D(n3630), .CP(
        n6091), .Q(mgmtsoc_master_rxtx_w[5]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[6]  ( .D(n3184), .CP(n6112), .Q(
        mgmtsoc_litespisdrphycore_source_payload_data[6]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[6]  ( .D(n3629), .CP(
        n6091), .Q(mgmtsoc_master_rxtx_w[6]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[6]  ( .D(N4249), .CP(n6054), .Q(
        interface3_bank_bus_dat_r[6]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[7]  ( .D(n3183), .CP(n6091), .Q(
        mgmtsoc_litespisdrphycore_source_payload_data[7]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[7]  ( .D(n3628), .CP(
        n6048), .Q(mgmtsoc_master_rxtx_w[7]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[7]  ( .D(N4250), .CP(n6043), .Q(
        interface3_bank_bus_dat_r[7]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[8]  ( .D(n3182), .CP(n6043), .Q(
        mgmtsoc_litespisdrphycore_source_payload_data[8]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[8]  ( .D(n3627), .CP(
        n6043), .Q(mgmtsoc_master_rxtx_w[8]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[8]  ( .D(N4251), .CP(n6043), .Q(
        interface3_bank_bus_dat_r[8]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[9]  ( .D(n3181), .CP(n6043), .Q(
        mgmtsoc_litespisdrphycore_source_payload_data[9]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[9]  ( .D(n3626), .CP(
        n6043), .Q(mgmtsoc_master_rxtx_w[9]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[10]  ( .D(n3180), .CP(n6043), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[10]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[10]  ( .D(n3625), 
        .CP(n6043), .Q(mgmtsoc_master_rxtx_w[10]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[11]  ( .D(n3179), .CP(n6089), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[11]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[11]  ( .D(n3624), 
        .CP(n6125), .Q(mgmtsoc_master_rxtx_w[11]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[11]  ( .D(N4254), .CP(n6101), .Q(
        interface3_bank_bus_dat_r[11]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[12]  ( .D(n3178), .CP(n6125), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[12]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[12]  ( .D(n3623), 
        .CP(n6100), .Q(mgmtsoc_master_rxtx_w[12]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[13]  ( .D(n3177), .CP(n6125), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[13]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[13]  ( .D(n3622), 
        .CP(n6026), .Q(mgmtsoc_master_rxtx_w[13]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[14]  ( .D(n3176), .CP(n6125), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[14]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[14]  ( .D(n3621), 
        .CP(n6044), .Q(mgmtsoc_master_rxtx_w[14]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[15]  ( .D(n3175), .CP(n6089), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[15]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[15]  ( .D(n3620), 
        .CP(n6044), .Q(mgmtsoc_master_rxtx_w[15]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[16]  ( .D(n3174), .CP(n6089), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[16]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[16]  ( .D(n3619), 
        .CP(n6044), .Q(mgmtsoc_master_rxtx_w[16]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[16]  ( .D(N4259), .CP(n6089), .Q(
        interface3_bank_bus_dat_r[16]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[17]  ( .D(n3173), .CP(n6044), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[17]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[17]  ( .D(n3618), 
        .CP(n6089), .Q(mgmtsoc_master_rxtx_w[17]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[18]  ( .D(n3172), .CP(n6045), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[18]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[18]  ( .D(n3617), 
        .CP(n6088), .Q(mgmtsoc_master_rxtx_w[18]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[19]  ( .D(n3171), .CP(n6045), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[19]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[19]  ( .D(n3616), 
        .CP(n6088), .Q(mgmtsoc_master_rxtx_w[19]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[20]  ( .D(n3170), .CP(n6045), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[20]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[20]  ( .D(n3615), 
        .CP(n6088), .Q(mgmtsoc_master_rxtx_w[20]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[21]  ( .D(n3169), .CP(n6045), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[21]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[21]  ( .D(n3614), 
        .CP(n6088), .Q(mgmtsoc_master_rxtx_w[21]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[22]  ( .D(n3168), .CP(n6048), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[22]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[22]  ( .D(n3613), 
        .CP(n6036), .Q(mgmtsoc_master_rxtx_w[22]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[23]  ( .D(n3167), .CP(n6041), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[23]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[23]  ( .D(n3612), 
        .CP(n6114), .Q(mgmtsoc_master_rxtx_w[23]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[24]  ( .D(n3166), .CP(n6036), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[24]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[24]  ( .D(n3611), 
        .CP(n6061), .Q(mgmtsoc_master_rxtx_w[24]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[24]  ( .D(N4267), .CP(n6059), .Q(
        interface3_bank_bus_dat_r[24]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[25]  ( .D(n3165), .CP(n6126), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[25]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[25]  ( .D(n3610), 
        .CP(n6022), .Q(mgmtsoc_master_rxtx_w[25]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[25]  ( .D(N4268), .CP(n6035), .Q(
        interface3_bank_bus_dat_r[25]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[26]  ( .D(n3164), .CP(n6034), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[26]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[26]  ( .D(n3609), 
        .CP(n6126), .Q(mgmtsoc_master_rxtx_w[26]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[26]  ( .D(N4269), .CP(n6035), .Q(
        interface3_bank_bus_dat_r[26]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[27]  ( .D(n3163), .CP(n6035), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[27]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[27]  ( .D(n3608), 
        .CP(n6035), .Q(mgmtsoc_master_rxtx_w[27]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[27]  ( .D(N4270), .CP(n6034), .Q(
        interface3_bank_bus_dat_r[27]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_in_reg[28]  ( .D(n3162), .CP(n6034), 
        .Q(mgmtsoc_litespisdrphycore_source_payload_data[28]) );
  dfnrq1 \mgmtsoc_master_rx_fifo_source_payload_data_reg[28]  ( .D(n3607), 
        .CP(n6034), .Q(mgmtsoc_master_rxtx_w[28]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[28]  ( .D(N4271), .CP(n6034), .Q(
        interface3_bank_bus_dat_r[28]) );
  dfnrq1 \dbg_uart_data_reg[4]  ( .D(n3279), .CP(n6034), .Q(
        dbg_uart_wishbone_dat_w[4]) );
  dfnrq1 \spi_master_mosi_storage_reg[4]  ( .D(n4541), .CP(n6034), .Q(
        spi_master_mosi[4]) );
  dfnrq1 \spi_master_mosi_data_reg[4]  ( .D(n3689), .CP(n6034), .Q(
        spi_master_mosi_data[4]) );
  dfnrq1 spi_mosi_reg ( .D(n3638), .CP(n6034), .Q(spi_mosi) );
  dfnrq1 \spi_master_miso_data_reg[0]  ( .D(n3704), .CP(n6035), .Q(
        spi_master_miso_data[0]) );
  dfnrq1 \spi_master_miso_data_reg[1]  ( .D(n3703), .CP(n6035), .Q(
        spi_master_miso_data[1]) );
  dfnrq1 \spi_master_miso_data_reg[2]  ( .D(n3702), .CP(n6035), .Q(
        spi_master_miso_data[2]) );
  dfnrq1 \spi_master_miso_data_reg[3]  ( .D(n3701), .CP(n6035), .Q(
        spi_master_miso_data[3]) );
  dfnrq1 \spi_master_miso_data_reg[4]  ( .D(n3700), .CP(n6035), .Q(
        spi_master_miso_data[4]) );
  dfnrq1 \spi_master_miso_data_reg[5]  ( .D(n3699), .CP(n6035), .Q(
        spi_master_miso_data[5]) );
  dfnrq1 \spi_master_miso_data_reg[6]  ( .D(n3698), .CP(n6035), .Q(
        spi_master_miso_data[6]) );
  dfnrq1 \spi_master_miso_data_reg[7]  ( .D(n3697), .CP(n6035), .Q(
        spi_master_miso_data[7]) );
  dfnrq1 \spi_master_miso_reg[7]  ( .D(n3639), .CP(n6035), .Q(
        spi_master_miso_status[7]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[7]  ( .D(N4592), .CP(n6034), .Q(
        interface9_bank_bus_dat_r[7]) );
  dfnrq1 \spi_master_miso_reg[6]  ( .D(n3640), .CP(n6034), .Q(
        spi_master_miso_status[6]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[6]  ( .D(N4591), .CP(n6126), .Q(
        interface9_bank_bus_dat_r[6]) );
  dfnrq1 \spi_master_miso_reg[5]  ( .D(n3641), .CP(n6034), .Q(
        spi_master_miso_status[5]) );
  dfnrq1 \spi_master_miso_reg[4]  ( .D(n3642), .CP(n6034), .Q(
        spi_master_miso_status[4]) );
  dfnrq1 \spi_master_miso_reg[3]  ( .D(n3643), .CP(n6126), .Q(
        spi_master_miso_status[3]) );
  dfnrq1 \spi_master_miso_reg[2]  ( .D(n3644), .CP(n6126), .Q(
        spi_master_miso_status[2]) );
  dfnrq1 \spi_master_miso_reg[1]  ( .D(n3645), .CP(n6126), .Q(
        spi_master_miso_status[1]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[1]  ( .D(N4586), .CP(n6035), .Q(
        interface9_bank_bus_dat_r[1]) );
  dfnrq1 \dbg_uart_data_reg[1]  ( .D(n3282), .CP(n6120), .Q(
        dbg_uart_wishbone_dat_w[1]) );
  dfnrq1 \spi_master_mosi_storage_reg[1]  ( .D(n4544), .CP(n6126), .Q(
        spi_master_mosi[1]) );
  dfnrq1 \spi_master_mosi_data_reg[1]  ( .D(n3692), .CP(n6035), .Q(
        spi_master_mosi_data[1]) );
  dfnrq1 \la_out_storage_reg[1]  ( .D(n4479), .CP(n6126), .Q(n133) );
  dfnrq1 \la_out_storage_reg[33]  ( .D(n4447), .CP(n6119), .Q(n101) );
  dfnrq1 \la_out_storage_reg[65]  ( .D(n4415), .CP(n6126), .Q(n69) );
  dfnrq1 \la_out_storage_reg[97]  ( .D(n4383), .CP(n6090), .Q(n37) );
  dfnrq1 \la_oe_storage_reg[1]  ( .D(n4351), .CP(n6100), .Q(csrbank6_oe0_w[1])
         );
  dfnrq1 \la_oe_storage_reg[33]  ( .D(n4319), .CP(n6090), .Q(csrbank6_oe1_w[1]) );
  dfnrq1 \la_oe_storage_reg[65]  ( .D(n4287), .CP(n6125), .Q(csrbank6_oe2_w[1]) );
  dfnrq1 \la_oe_storage_reg[97]  ( .D(n4255), .CP(n6090), .Q(csrbank6_oe3_w[1]) );
  dfnrq1 \la_ien_storage_reg[1]  ( .D(n4223), .CP(n6090), .Q(
        csrbank6_ien0_w[1]) );
  dfnrq1 \la_ien_storage_reg[33]  ( .D(n4191), .CP(n6090), .Q(
        csrbank6_ien1_w[1]) );
  dfnrq1 \la_ien_storage_reg[65]  ( .D(n4159), .CP(n6090), .Q(
        csrbank6_ien2_w[1]) );
  dfnrq1 \la_ien_storage_reg[97]  ( .D(n4127), .CP(n6039), .Q(
        csrbank6_ien3_w[1]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[1]  ( .D(N4464), .CP(n6048), .Q(
        interface6_bank_bus_dat_r[1]) );
  dfnrq1 \storage_reg[15][1]  ( .D(n4038), .CP(n6036), .Q(\storage[15][1] ) );
  dfnrq1 \storage_reg[14][1]  ( .D(n4030), .CP(n6041), .Q(\storage[14][1] ) );
  dfnrq1 \storage_reg[13][1]  ( .D(n4022), .CP(n6038), .Q(\storage[13][1] ) );
  dfnrq1 \storage_reg[12][1]  ( .D(n4014), .CP(n6041), .Q(\storage[12][1] ) );
  dfnrq1 \storage_reg[11][1]  ( .D(n4006), .CP(n6040), .Q(\storage[11][1] ) );
  dfnrq1 \storage_reg[10][1]  ( .D(n3998), .CP(n6095), .Q(\storage[10][1] ) );
  dfnrq1 \storage_reg[9][1]  ( .D(n3990), .CP(n6036), .Q(\storage[9][1] ) );
  dfnrq1 \storage_reg[8][1]  ( .D(n3982), .CP(n6036), .Q(\storage[8][1] ) );
  dfnrq1 \storage_reg[7][1]  ( .D(n3974), .CP(n6036), .Q(\storage[7][1] ) );
  dfnrq1 \storage_reg[6][1]  ( .D(n3966), .CP(n6036), .Q(\storage[6][1] ) );
  dfnrq1 \storage_reg[5][1]  ( .D(n3958), .CP(n6036), .Q(\storage[5][1] ) );
  dfnrq1 \storage_reg[4][1]  ( .D(n3950), .CP(n6036), .Q(\storage[4][1] ) );
  dfnrq1 \storage_reg[3][1]  ( .D(n3942), .CP(n6036), .Q(\storage[3][1] ) );
  dfnrq1 \storage_reg[2][1]  ( .D(n3934), .CP(n6039), .Q(\storage[2][1] ) );
  dfnrq1 \storage_reg[1][1]  ( .D(n3926), .CP(n6048), .Q(\storage[1][1] ) );
  dfnrq1 \storage_reg[0][1]  ( .D(n3918), .CP(n6036), .Q(\storage[0][1] ) );
  dfnrq1 \memdat_1_reg[1]  ( .D(n3892), .CP(n6041), .Q(
        uart_tx_fifo_fifo_out_payload_data[1]) );
  dfnrq1 \spimaster_storage_reg[1]  ( .D(n3719), .CP(n6114), .Q(
        spi_master_clk_divider0[1]) );
  dfnrq1 \spi_master_cs_storage_reg[1]  ( .D(n3680), .CP(n6039), .Q(
        csrbank9_cs0_w[1]) );
  dfnrq1 \spi_master_control_storage_reg[1]  ( .D(n3661), .CP(n6041), .Q(
        csrbank9_control0_w[1]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[1]  ( .D(n3601), .CP(
        n6039), .Q(mgmtsoc_port_master_user_port_sink_payload_data[1]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[1]  ( .D(n3558), .CP(n6037), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_len[1]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_len_reg[1]  ( .D(n3569), .CP(
        n6037), .Q(mgmtsoc_port_master_user_port_sink_payload_len[1]) );
  dfnrq1 \mgmtsoc_litespimmap_storage_reg[1]  ( .D(n3533), .CP(n6037), .Q(
        mgmtsoc_litespimmap_spi_dummy_bits[1]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[1]  ( .D(N4244), .CP(n6037), .Q(
        interface3_bank_bus_dat_r[1]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_storage_reg[1]  ( .D(n3510), .CP(n6037), 
        .Q(mgmtsoc_litespisdrphycore_div[1]) );
  dfnrq1 \interface4_bank_bus_dat_r_reg[1]  ( .D(N4293), .CP(n6037), .Q(
        interface4_bank_bus_dat_r[1]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[1]  ( .D(n3465), .CP(n6037), .Q(
        csrbank10_reload0_w[1]) );
  dfnrq1 \mgmtsoc_load_storage_reg[1]  ( .D(n3433), .CP(n6037), .Q(
        csrbank10_load0_w[1]) );
  dfnrq1 \mgmtsoc_value_reg[1]  ( .D(N5401), .CP(n6114), .Q(mgmtsoc_value[1])
         );
  dfnrq1 \mgmtsoc_value_status_reg[1]  ( .D(n3499), .CP(n6047), .Q(
        csrbank10_value_w[1]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[1]  ( .D(N4695), .CP(n6038), .Q(
        interface10_bank_bus_dat_r[1]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[1]  ( .D(n3326), .CP(n6036), .Q(
        csrbank0_scratch0_w[1]) );
  dfnrq1 \user_irq_ena_storage_reg[1]  ( .D(n4483), .CP(n6037), .Q(n6132) );
  dfnrq1 \interface19_bank_bus_dat_r_reg[1]  ( .D(N4996), .CP(n6114), .Q(
        interface19_bank_bus_dat_r[1]) );
  dfnrq1 \uart_enable_storage_reg[1]  ( .D(n3909), .CP(n6047), .Q(
        csrbank11_ev_enable0_w[1]) );
  dfnrq1 \uart_pending_r_reg[1]  ( .D(n3907), .CP(n6038), .Q(uart_pending_r[1]) );
  dfnrq1 \uart_rx_fifo_consume_reg[0]  ( .D(n4066), .CP(n6038), .Q(
        uart_rx_fifo_rdport_adr[0]) );
  dfnrq1 \uart_rx_fifo_consume_reg[1]  ( .D(n4065), .CP(n6038), .Q(
        uart_rx_fifo_rdport_adr[1]) );
  dfnrq1 \uart_rx_fifo_consume_reg[2]  ( .D(n4064), .CP(n6038), .Q(
        uart_rx_fifo_rdport_adr[2]) );
  dfnrq1 \uart_rx_fifo_consume_reg[3]  ( .D(n4063), .CP(n6038), .Q(
        uart_rx_fifo_rdport_adr[3]) );
  dfnrq1 \uart_rx_fifo_level0_reg[1]  ( .D(n4054), .CP(n6038), .Q(
        uart_rx_fifo_level0[1]) );
  dfnrq1 \uart_rx_fifo_level0_reg[0]  ( .D(n4058), .CP(n6038), .Q(
        uart_rx_fifo_level0[0]) );
  dfnrq1 \uart_rx_fifo_level0_reg[4]  ( .D(n4057), .CP(n6038), .Q(
        uart_rx_fifo_level0[4]) );
  dfnrq1 \uart_rx_fifo_level0_reg[3]  ( .D(n4056), .CP(n6038), .Q(
        uart_rx_fifo_level0[3]) );
  dfnrq1 \uart_rx_fifo_level0_reg[2]  ( .D(n4055), .CP(n6039), .Q(
        uart_rx_fifo_level0[2]) );
  dfnrq1 \uart_rx_fifo_produce_reg[0]  ( .D(n4062), .CP(n6039), .Q(
        uart_rx_fifo_produce[0]) );
  dfnrq1 \uart_rx_fifo_produce_reg[1]  ( .D(n4061), .CP(n6039), .Q(
        uart_rx_fifo_produce[1]) );
  dfnrq1 \uart_rx_fifo_produce_reg[2]  ( .D(n4060), .CP(n6039), .Q(
        uart_rx_fifo_produce[2]) );
  dfnrq1 \uart_rx_fifo_produce_reg[3]  ( .D(n4059), .CP(n6039), .Q(
        uart_rx_fifo_produce[3]) );
  dfnrq1 \storage_1_reg[15][0]  ( .D(n3864), .CP(n6039), .Q(\storage_1[15][0] ) );
  dfnrq1 \storage_1_reg[15][1]  ( .D(n3863), .CP(n6039), .Q(\storage_1[15][1] ) );
  dfnrq1 \storage_1_reg[15][2]  ( .D(n3862), .CP(n6039), .Q(\storage_1[15][2] ) );
  dfnrq1 \storage_1_reg[15][3]  ( .D(n3861), .CP(n6113), .Q(\storage_1[15][3] ) );
  dfnrq1 \storage_1_reg[15][4]  ( .D(n3860), .CP(n6049), .Q(\storage_1[15][4] ) );
  dfnrq1 \storage_1_reg[15][5]  ( .D(n3859), .CP(n6087), .Q(\storage_1[15][5] ) );
  dfnrq1 \storage_1_reg[15][6]  ( .D(n3858), .CP(n6042), .Q(\storage_1[15][6] ) );
  dfnrq1 \storage_1_reg[15][7]  ( .D(n3857), .CP(n6043), .Q(\storage_1[15][7] ) );
  dfnrq1 \storage_1_reg[13][0]  ( .D(n3848), .CP(n6049), .Q(\storage_1[13][0] ) );
  dfnrq1 \storage_1_reg[13][1]  ( .D(n3847), .CP(n6087), .Q(\storage_1[13][1] ) );
  dfnrq1 \storage_1_reg[13][2]  ( .D(n3846), .CP(n6113), .Q(\storage_1[13][2] ) );
  dfnrq1 \storage_1_reg[13][3]  ( .D(n3845), .CP(n6087), .Q(\storage_1[13][3] ) );
  dfnrq1 \storage_1_reg[13][4]  ( .D(n3844), .CP(n6043), .Q(\storage_1[13][4] ) );
  dfnrq1 \storage_1_reg[13][5]  ( .D(n3843), .CP(n6040), .Q(\storage_1[13][5] ) );
  dfnrq1 \storage_1_reg[13][6]  ( .D(n3842), .CP(n6042), .Q(\storage_1[13][6] ) );
  dfnrq1 \storage_1_reg[13][7]  ( .D(n3841), .CP(n6043), .Q(\storage_1[13][7] ) );
  dfnrq1 \storage_1_reg[11][0]  ( .D(n3832), .CP(n6047), .Q(\storage_1[11][0] ) );
  dfnrq1 \storage_1_reg[11][1]  ( .D(n3831), .CP(n6098), .Q(\storage_1[11][1] ) );
  dfnrq1 \storage_1_reg[11][2]  ( .D(n3830), .CP(n6097), .Q(\storage_1[11][2] ) );
  dfnrq1 \storage_1_reg[11][3]  ( .D(n3829), .CP(n6026), .Q(\storage_1[11][3] ) );
  dfnrq1 \storage_1_reg[11][4]  ( .D(n3828), .CP(n6084), .Q(\storage_1[11][4] ) );
  dfnrq1 \storage_1_reg[11][5]  ( .D(n3827), .CP(n6092), .Q(\storage_1[11][5] ) );
  dfnrq1 \storage_1_reg[11][6]  ( .D(n3826), .CP(n6102), .Q(\storage_1[11][6] ) );
  dfnrq1 \storage_1_reg[11][7]  ( .D(n3825), .CP(n6093), .Q(\storage_1[11][7] ) );
  dfnrq1 \storage_1_reg[9][0]  ( .D(n3816), .CP(n6095), .Q(\storage_1[9][0] )
         );
  dfnrq1 \storage_1_reg[9][1]  ( .D(n3815), .CP(n6077), .Q(\storage_1[9][1] )
         );
  dfnrq1 \storage_1_reg[9][2]  ( .D(n3814), .CP(n6083), .Q(\storage_1[9][2] )
         );
  dfnrq1 \storage_1_reg[9][3]  ( .D(n3813), .CP(n6082), .Q(\storage_1[9][3] )
         );
  dfnrq1 \storage_1_reg[9][4]  ( .D(n3812), .CP(n6124), .Q(\storage_1[9][4] )
         );
  dfnrq1 \storage_1_reg[9][5]  ( .D(n3811), .CP(n6095), .Q(\storage_1[9][5] )
         );
  dfnrq1 \storage_1_reg[9][6]  ( .D(n3810), .CP(n6124), .Q(\storage_1[9][6] )
         );
  dfnrq1 \storage_1_reg[9][7]  ( .D(n3809), .CP(n6092), .Q(\storage_1[9][7] )
         );
  dfnrq1 \storage_1_reg[7][0]  ( .D(n3800), .CP(n6124), .Q(\storage_1[7][0] )
         );
  dfnrq1 \storage_1_reg[7][1]  ( .D(n3799), .CP(n6124), .Q(\storage_1[7][1] )
         );
  dfnrq1 \storage_1_reg[7][2]  ( .D(n3798), .CP(n6092), .Q(\storage_1[7][2] )
         );
  dfnrq1 \storage_1_reg[7][3]  ( .D(n3797), .CP(n6102), .Q(\storage_1[7][3] )
         );
  dfnrq1 \storage_1_reg[7][4]  ( .D(n3796), .CP(n6094), .Q(\storage_1[7][4] )
         );
  dfnrq1 \storage_1_reg[7][5]  ( .D(n3795), .CP(n6094), .Q(\storage_1[7][5] )
         );
  dfnrq1 \storage_1_reg[7][6]  ( .D(n3794), .CP(n6094), .Q(\storage_1[7][6] )
         );
  dfnrq1 \storage_1_reg[7][7]  ( .D(n3793), .CP(n6094), .Q(\storage_1[7][7] )
         );
  dfnrq1 \storage_1_reg[5][0]  ( .D(n3784), .CP(n6094), .Q(\storage_1[5][0] )
         );
  dfnrq1 \storage_1_reg[5][1]  ( .D(n3783), .CP(n6094), .Q(\storage_1[5][1] )
         );
  dfnrq1 \storage_1_reg[5][2]  ( .D(n3782), .CP(n6094), .Q(\storage_1[5][2] )
         );
  dfnrq1 \storage_1_reg[5][3]  ( .D(n3781), .CP(n6094), .Q(\storage_1[5][3] )
         );
  dfnrq1 \storage_1_reg[5][4]  ( .D(n3780), .CP(n6095), .Q(\storage_1[5][4] )
         );
  dfnrq1 \storage_1_reg[5][5]  ( .D(n3779), .CP(n6095), .Q(\storage_1[5][5] )
         );
  dfnrq1 \storage_1_reg[5][6]  ( .D(n3778), .CP(n6095), .Q(\storage_1[5][6] )
         );
  dfnrq1 \storage_1_reg[5][7]  ( .D(n3777), .CP(n6095), .Q(\storage_1[5][7] )
         );
  dfnrq1 \storage_1_reg[3][0]  ( .D(n3768), .CP(n6095), .Q(\storage_1[3][0] )
         );
  dfnrq1 \storage_1_reg[3][1]  ( .D(n3767), .CP(n6095), .Q(\storage_1[3][1] )
         );
  dfnrq1 \storage_1_reg[3][2]  ( .D(n3766), .CP(n6095), .Q(\storage_1[3][2] )
         );
  dfnrq1 \storage_1_reg[3][3]  ( .D(n3765), .CP(n6095), .Q(\storage_1[3][3] )
         );
  dfnrq1 \storage_1_reg[3][4]  ( .D(n3764), .CP(n6083), .Q(\storage_1[3][4] )
         );
  dfnrq1 \storage_1_reg[3][5]  ( .D(n3763), .CP(n6122), .Q(\storage_1[3][5] )
         );
  dfnrq1 \storage_1_reg[3][6]  ( .D(n3762), .CP(n6083), .Q(\storage_1[3][6] )
         );
  dfnrq1 \storage_1_reg[3][7]  ( .D(n3761), .CP(n6122), .Q(\storage_1[3][7] )
         );
  dfnrq1 \storage_1_reg[1][0]  ( .D(n3752), .CP(n6083), .Q(\storage_1[1][0] )
         );
  dfnrq1 \storage_1_reg[1][1]  ( .D(n3751), .CP(n6083), .Q(\storage_1[1][1] )
         );
  dfnrq1 \storage_1_reg[1][2]  ( .D(n3750), .CP(n6083), .Q(\storage_1[1][2] )
         );
  dfnrq1 \storage_1_reg[1][3]  ( .D(n3749), .CP(n6083), .Q(\storage_1[1][3] )
         );
  dfnrq1 \storage_1_reg[1][4]  ( .D(n3748), .CP(n6096), .Q(\storage_1[1][4] )
         );
  dfnrq1 \storage_1_reg[1][5]  ( .D(n3747), .CP(n6096), .Q(\storage_1[1][5] )
         );
  dfnrq1 \storage_1_reg[1][6]  ( .D(n3746), .CP(n6096), .Q(\storage_1[1][6] )
         );
  dfnrq1 \storage_1_reg[1][7]  ( .D(n3745), .CP(n6096), .Q(\storage_1[1][7] )
         );
  dfnrq1 \storage_1_reg[14][0]  ( .D(n3856), .CP(n6096), .Q(\storage_1[14][0] ) );
  dfnrq1 \storage_1_reg[14][1]  ( .D(n3855), .CP(n6096), .Q(\storage_1[14][1] ) );
  dfnrq1 \storage_1_reg[14][2]  ( .D(n3854), .CP(n6096), .Q(\storage_1[14][2] ) );
  dfnrq1 \storage_1_reg[14][3]  ( .D(n3853), .CP(n6096), .Q(\storage_1[14][3] ) );
  dfnrq1 \storage_1_reg[14][4]  ( .D(n3852), .CP(n6084), .Q(\storage_1[14][4] ) );
  dfnrq1 \storage_1_reg[14][5]  ( .D(n3851), .CP(n6123), .Q(\storage_1[14][5] ) );
  dfnrq1 \storage_1_reg[14][6]  ( .D(n3850), .CP(n6095), .Q(\storage_1[14][6] ) );
  dfnrq1 \storage_1_reg[14][7]  ( .D(n3849), .CP(n6123), .Q(\storage_1[14][7] ) );
  dfnrq1 \storage_1_reg[12][0]  ( .D(n3840), .CP(n6123), .Q(\storage_1[12][0] ) );
  dfnrq1 \storage_1_reg[12][1]  ( .D(n3839), .CP(n6123), .Q(\storage_1[12][1] ) );
  dfnrq1 \storage_1_reg[12][2]  ( .D(n3838), .CP(n6124), .Q(\storage_1[12][2] ) );
  dfnrq1 \storage_1_reg[12][3]  ( .D(n3837), .CP(n6123), .Q(\storage_1[12][3] ) );
  dfnrq1 \storage_1_reg[12][4]  ( .D(n3836), .CP(n6076), .Q(\storage_1[12][4] ) );
  dfnrq1 \storage_1_reg[12][5]  ( .D(n3835), .CP(n6076), .Q(\storage_1[12][5] ) );
  dfnrq1 \storage_1_reg[12][6]  ( .D(n3834), .CP(n6097), .Q(\storage_1[12][6] ) );
  dfnrq1 \storage_1_reg[12][7]  ( .D(n3833), .CP(n6076), .Q(\storage_1[12][7] ) );
  dfnrq1 \storage_1_reg[10][0]  ( .D(n3824), .CP(n6097), .Q(\storage_1[10][0] ) );
  dfnrq1 \storage_1_reg[10][1]  ( .D(n3823), .CP(n6097), .Q(\storage_1[10][1] ) );
  dfnrq1 \storage_1_reg[10][2]  ( .D(n3822), .CP(n6097), .Q(\storage_1[10][2] ) );
  dfnrq1 \storage_1_reg[10][3]  ( .D(n3821), .CP(n6051), .Q(\storage_1[10][3] ) );
  dfnrq1 \storage_1_reg[10][4]  ( .D(n3820), .CP(n6032), .Q(\storage_1[10][4] ) );
  dfnrq1 \storage_1_reg[10][5]  ( .D(n3819), .CP(n6032), .Q(\storage_1[10][5] ) );
  dfnrq1 \storage_1_reg[10][6]  ( .D(n3818), .CP(n6098), .Q(\storage_1[10][6] ) );
  dfnrq1 \storage_1_reg[10][7]  ( .D(n3817), .CP(n6022), .Q(\storage_1[10][7] ) );
  dfnrq1 \storage_1_reg[8][0]  ( .D(n3808), .CP(n6051), .Q(\storage_1[8][0] )
         );
  dfnrq1 \storage_1_reg[8][1]  ( .D(n3807), .CP(n6032), .Q(\storage_1[8][1] )
         );
  dfnrq1 \storage_1_reg[8][2]  ( .D(n3806), .CP(n6022), .Q(\storage_1[8][2] )
         );
  dfnrq1 \storage_1_reg[8][3]  ( .D(n3805), .CP(n6088), .Q(\storage_1[8][3] )
         );
  dfnrq1 \storage_1_reg[8][4]  ( .D(n3804), .CP(n6125), .Q(\storage_1[8][4] )
         );
  dfnrq1 \storage_1_reg[8][5]  ( .D(n3803), .CP(n6100), .Q(\storage_1[8][5] )
         );
  dfnrq1 \storage_1_reg[8][6]  ( .D(n3802), .CP(n6045), .Q(\storage_1[8][6] )
         );
  dfnrq1 \storage_1_reg[8][7]  ( .D(n3801), .CP(n6044), .Q(\storage_1[8][7] )
         );
  dfnrq1 \storage_1_reg[6][0]  ( .D(n3792), .CP(n6091), .Q(\storage_1[6][0] )
         );
  dfnrq1 \storage_1_reg[6][1]  ( .D(n3791), .CP(n6039), .Q(\storage_1[6][1] )
         );
  dfnrq1 \storage_1_reg[6][2]  ( .D(n3790), .CP(n6026), .Q(\storage_1[6][2] )
         );
  dfnrq1 \storage_1_reg[6][3]  ( .D(n3789), .CP(n6094), .Q(\storage_1[6][3] )
         );
  dfnrq1 \storage_1_reg[6][4]  ( .D(n3788), .CP(n6101), .Q(\storage_1[6][4] )
         );
  dfnrq1 \storage_1_reg[6][5]  ( .D(n3787), .CP(n6059), .Q(\storage_1[6][5] )
         );
  dfnrq1 \storage_1_reg[6][6]  ( .D(n3786), .CP(n6125), .Q(\storage_1[6][6] )
         );
  dfnrq1 \storage_1_reg[6][7]  ( .D(n3785), .CP(n6101), .Q(\storage_1[6][7] )
         );
  dfnrq1 \storage_1_reg[4][0]  ( .D(n3776), .CP(n6100), .Q(\storage_1[4][0] )
         );
  dfnrq1 \storage_1_reg[4][1]  ( .D(n3775), .CP(n6026), .Q(\storage_1[4][1] )
         );
  dfnrq1 \storage_1_reg[4][2]  ( .D(n3774), .CP(n6029), .Q(\storage_1[4][2] )
         );
  dfnrq1 \storage_1_reg[4][3]  ( .D(n3773), .CP(n6094), .Q(\storage_1[4][3] )
         );
  dfnrq1 \storage_1_reg[4][4]  ( .D(n3772), .CP(n6101), .Q(\storage_1[4][4] )
         );
  dfnrq1 \storage_1_reg[4][5]  ( .D(n3771), .CP(n6100), .Q(\storage_1[4][5] )
         );
  dfnrq1 \storage_1_reg[4][6]  ( .D(n3770), .CP(n6125), .Q(\storage_1[4][6] )
         );
  dfnrq1 \storage_1_reg[4][7]  ( .D(n3769), .CP(n6026), .Q(\storage_1[4][7] )
         );
  dfnrq1 \storage_1_reg[2][0]  ( .D(n3760), .CP(n6029), .Q(\storage_1[2][0] )
         );
  dfnrq1 \storage_1_reg[2][1]  ( .D(n3759), .CP(n6094), .Q(\storage_1[2][1] )
         );
  dfnrq1 \storage_1_reg[2][2]  ( .D(n3758), .CP(n6024), .Q(\storage_1[2][2] )
         );
  dfnrq1 \storage_1_reg[2][3]  ( .D(n3757), .CP(n6026), .Q(\storage_1[2][3] )
         );
  dfnrq1 \storage_1_reg[2][4]  ( .D(n3756), .CP(n6029), .Q(\storage_1[2][4] )
         );
  dfnrq1 \storage_1_reg[2][5]  ( .D(n3755), .CP(n6057), .Q(\storage_1[2][5] )
         );
  dfnrq1 \storage_1_reg[2][6]  ( .D(n3754), .CP(n6112), .Q(\storage_1[2][6] )
         );
  dfnrq1 \storage_1_reg[2][7]  ( .D(n3753), .CP(n6094), .Q(\storage_1[2][7] )
         );
  dfnrq1 \storage_1_reg[0][0]  ( .D(n3744), .CP(n6088), .Q(\storage_1[0][0] )
         );
  dfnrq1 \storage_1_reg[0][1]  ( .D(n3743), .CP(n6061), .Q(\storage_1[0][1] )
         );
  dfnrq1 \storage_1_reg[0][2]  ( .D(n3741), .CP(n6041), .Q(\storage_1[0][2] )
         );
  dfnrq1 \storage_1_reg[0][3]  ( .D(n3739), .CP(n6097), .Q(\storage_1[0][3] )
         );
  dfnrq1 \storage_1_reg[0][4]  ( .D(n3737), .CP(n6097), .Q(\storage_1[0][4] )
         );
  dfnrq1 \storage_1_reg[0][5]  ( .D(n3735), .CP(n6097), .Q(\storage_1[0][5] )
         );
  dfnrq1 \storage_1_reg[0][6]  ( .D(n3733), .CP(n6097), .Q(\storage_1[0][6] )
         );
  dfnrq1 \storage_1_reg[0][7]  ( .D(n3731), .CP(n6097), .Q(\storage_1[0][7] )
         );
  dfnrq1 uart_rx_fifo_readable_reg ( .D(n4053), .CP(n6097), .Q(
        \uart_status_status[1] ) );
  dfnrq1 uart_rx_trigger_d_reg ( .D(N5710), .CP(n6097), .Q(uart_rx_trigger_d)
         );
  dfnrq1 uart_rx_pending_reg ( .D(n3906), .CP(n6097), .Q(
        uart_pending_status[1]) );
  dfnrq1 \memdat_3_reg[1]  ( .D(n3742), .CP(n6098), .Q(
        uart_rx_fifo_fifo_out_payload_data[1]) );
  dfnrq1 \interface11_bank_bus_dat_r_reg[1]  ( .D(N4773), .CP(n6098), .Q(
        interface11_bank_bus_dat_r[1]) );
  dfnrq1 \memdat_3_reg[2]  ( .D(n3740), .CP(n6098), .Q(
        uart_rx_fifo_fifo_out_payload_data[2]) );
  dfnrq1 \interface11_bank_bus_dat_r_reg[2]  ( .D(N4774), .CP(n6098), .Q(
        interface11_bank_bus_dat_r[2]) );
  dfnrq1 \dbg_uart_data_reg[2]  ( .D(n3281), .CP(n6098), .Q(
        dbg_uart_wishbone_dat_w[2]) );
  dfnrq1 \spi_master_mosi_storage_reg[2]  ( .D(n4543), .CP(n6088), .Q(
        spi_master_mosi[2]) );
  dfnrq1 \spi_master_mosi_data_reg[2]  ( .D(n3691), .CP(n6077), .Q(
        spi_master_mosi_data[2]) );
  dfnrq1 \user_irq_ena_storage_reg[2]  ( .D(n4482), .CP(n6121), .Q(n6131) );
  dfnrq1 \interface19_bank_bus_dat_r_reg[2]  ( .D(N4997), .CP(n6077), .Q(
        interface19_bank_bus_dat_r[2]) );
  dfnrq1 \la_out_storage_reg[2]  ( .D(n4478), .CP(n6121), .Q(n132) );
  dfnrq1 \la_out_storage_reg[34]  ( .D(n4446), .CP(n6077), .Q(n100) );
  dfnrq1 \la_out_storage_reg[66]  ( .D(n4414), .CP(n6077), .Q(n68) );
  dfnrq1 \la_out_storage_reg[98]  ( .D(n4382), .CP(n6077), .Q(n36) );
  dfnrq1 \la_oe_storage_reg[2]  ( .D(n4350), .CP(n6077), .Q(csrbank6_oe0_w[2])
         );
  dfnrq1 \la_oe_storage_reg[34]  ( .D(n4318), .CP(n6091), .Q(csrbank6_oe1_w[2]) );
  dfnrq1 \la_oe_storage_reg[66]  ( .D(n4286), .CP(n6101), .Q(csrbank6_oe2_w[2]) );
  dfnrq1 \la_oe_storage_reg[98]  ( .D(n4254), .CP(n6087), .Q(csrbank6_oe3_w[2]) );
  dfnrq1 \la_ien_storage_reg[2]  ( .D(n4222), .CP(n6094), .Q(
        csrbank6_ien0_w[2]) );
  dfnrq1 \la_ien_storage_reg[34]  ( .D(n4190), .CP(n6029), .Q(
        csrbank6_ien1_w[2]) );
  dfnrq1 \la_ien_storage_reg[66]  ( .D(n4158), .CP(n6091), .Q(
        csrbank6_ien2_w[2]) );
  dfnrq1 \la_ien_storage_reg[98]  ( .D(n4126), .CP(n6093), .Q(
        csrbank6_ien3_w[2]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[2]  ( .D(N4465), .CP(n6078), .Q(
        interface6_bank_bus_dat_r[2]) );
  dfnrq1 \storage_reg[15][2]  ( .D(n4037), .CP(n6087), .Q(\storage[15][2] ) );
  dfnrq1 \storage_reg[14][2]  ( .D(n4029), .CP(n6087), .Q(\storage[14][2] ) );
  dfnrq1 \storage_reg[13][2]  ( .D(n4021), .CP(n6087), .Q(\storage[13][2] ) );
  dfnrq1 \storage_reg[12][2]  ( .D(n4013), .CP(n6087), .Q(\storage[12][2] ) );
  dfnrq1 \storage_reg[11][2]  ( .D(n4005), .CP(n6087), .Q(\storage[11][2] ) );
  dfnrq1 \storage_reg[10][2]  ( .D(n3997), .CP(n6087), .Q(\storage[10][2] ) );
  dfnrq1 \storage_reg[9][2]  ( .D(n3989), .CP(n6087), .Q(\storage[9][2] ) );
  dfnrq1 \storage_reg[8][2]  ( .D(n3981), .CP(n6087), .Q(\storage[8][2] ) );
  dfnrq1 \storage_reg[7][2]  ( .D(n3973), .CP(n6125), .Q(\storage[7][2] ) );
  dfnrq1 \storage_reg[6][2]  ( .D(n3965), .CP(n6045), .Q(\storage[6][2] ) );
  dfnrq1 \storage_reg[5][2]  ( .D(n3957), .CP(n6091), .Q(\storage[5][2] ) );
  dfnrq1 \storage_reg[4][2]  ( .D(n3949), .CP(n6039), .Q(\storage[4][2] ) );
  dfnrq1 \storage_reg[3][2]  ( .D(n3941), .CP(n6026), .Q(\storage[3][2] ) );
  dfnrq1 \storage_reg[2][2]  ( .D(n3933), .CP(n6029), .Q(\storage[2][2] ) );
  dfnrq1 \storage_reg[1][2]  ( .D(n3925), .CP(n6057), .Q(\storage[1][2] ) );
  dfnrq1 \storage_reg[0][2]  ( .D(n3917), .CP(n6094), .Q(\storage[0][2] ) );
  dfnrq1 \memdat_1_reg[2]  ( .D(n3893), .CP(n6091), .Q(
        uart_tx_fifo_fifo_out_payload_data[2]) );
  dfnrq1 \spi_master_cs_storage_reg[2]  ( .D(n3679), .CP(n6091), .Q(
        csrbank9_cs0_w[2]) );
  dfnrq1 \spi_master_control_storage_reg[2]  ( .D(n3660), .CP(n6091), .Q(
        csrbank9_control0_w[2]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[2]  ( .D(N4587), .CP(n6091), .Q(
        interface9_bank_bus_dat_r[2]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[2]  ( .D(n3600), .CP(
        n6091), .Q(mgmtsoc_port_master_user_port_sink_payload_data[2]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[2]  ( .D(n3557), .CP(n6091), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_len[2]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_len_reg[2]  ( .D(n3568), .CP(
        n6091), .Q(mgmtsoc_port_master_user_port_sink_payload_len[2]) );
  dfnrq1 \mgmtsoc_litespimmap_storage_reg[2]  ( .D(n3532), .CP(n6091), .Q(
        mgmtsoc_litespimmap_spi_dummy_bits[2]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[2]  ( .D(N4245), .CP(n6090), .Q(
        interface3_bank_bus_dat_r[2]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_storage_reg[2]  ( .D(n3509), .CP(n6090), 
        .Q(mgmtsoc_litespisdrphycore_div[2]) );
  dfnrq1 \interface4_bank_bus_dat_r_reg[2]  ( .D(N4294), .CP(n6090), .Q(
        interface4_bank_bus_dat_r[2]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[2]  ( .D(n3464), .CP(n6090), .Q(
        csrbank10_reload0_w[2]) );
  dfnrq1 \mgmtsoc_load_storage_reg[2]  ( .D(n3432), .CP(n6090), .Q(
        csrbank10_load0_w[2]) );
  dfnrq1 \mgmtsoc_value_reg[2]  ( .D(N5402), .CP(n6090), .Q(mgmtsoc_value[2])
         );
  dfnrq1 \mgmtsoc_value_status_reg[2]  ( .D(n3498), .CP(n6090), .Q(
        csrbank10_value_w[2]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[2]  ( .D(N4696), .CP(n6090), .Q(
        interface10_bank_bus_dat_r[2]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[2]  ( .D(n3325), .CP(n6089), .Q(
        csrbank0_scratch0_w[2]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[2]  ( .D(N4101), .CP(n6089), .Q(
        interface0_bank_bus_dat_r[2]) );
  dfnrq1 \dbg_uart_data_reg[10]  ( .D(n3273), .CP(n6089), .Q(
        dbg_uart_wishbone_dat_w[10]) );
  dfnrq1 \la_out_storage_reg[10]  ( .D(n4470), .CP(n6089), .Q(n124) );
  dfnrq1 \la_out_storage_reg[42]  ( .D(n4438), .CP(n6089), .Q(n92) );
  dfnrq1 \la_out_storage_reg[74]  ( .D(n4406), .CP(n6089), .Q(n60) );
  dfnrq1 \la_out_storage_reg[106]  ( .D(n4374), .CP(n6089), .Q(n28) );
  dfnrq1 \la_oe_storage_reg[10]  ( .D(n4342), .CP(n6089), .Q(
        csrbank6_oe0_w[10]) );
  dfnrq1 \la_oe_storage_reg[42]  ( .D(n4310), .CP(n6088), .Q(
        csrbank6_oe1_w[10]) );
  dfnrq1 \la_oe_storage_reg[74]  ( .D(n4278), .CP(n6088), .Q(
        csrbank6_oe2_w[10]) );
  dfnrq1 \la_oe_storage_reg[106]  ( .D(n4246), .CP(n6088), .Q(
        csrbank6_oe3_w[10]) );
  dfnrq1 \la_ien_storage_reg[10]  ( .D(n4214), .CP(n6088), .Q(
        csrbank6_ien0_w[10]) );
  dfnrq1 \la_ien_storage_reg[42]  ( .D(n4182), .CP(n6088), .Q(
        csrbank6_ien1_w[10]) );
  dfnrq1 \la_ien_storage_reg[74]  ( .D(n4150), .CP(n6088), .Q(
        csrbank6_ien2_w[10]) );
  dfnrq1 \la_ien_storage_reg[106]  ( .D(n4118), .CP(n6093), .Q(
        csrbank6_ien3_w[10]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[10]  ( .D(N4473), .CP(n6095), .Q(
        interface6_bank_bus_dat_r[10]) );
  dfnrq1 \spimaster_storage_reg[10]  ( .D(n3710), .CP(n6084), .Q(
        spi_master_clk_divider0[10]) );
  dfnrq1 \spi_master_cs_storage_reg[10]  ( .D(n3671), .CP(n6092), .Q(
        csrbank9_cs0_w[10]) );
  dfnrq1 \spi_master_control_storage_reg[10]  ( .D(n3652), .CP(n6093), .Q(
        spi_master_length0[2]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[10]  ( .D(N4595), .CP(n6092), .Q(
        interface9_bank_bus_dat_r[10]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[10]  ( .D(n3592), 
        .CP(n6102), .Q(mgmtsoc_port_master_user_port_sink_payload_data[10]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[10]  ( .D(n3549), .CP(n6093), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_width[2]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[10]  ( .D(N4253), .CP(n6096), .Q(
        interface3_bank_bus_dat_r[10]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[10]  ( .D(n3456), .CP(n6095), .Q(
        csrbank10_reload0_w[10]) );
  dfnrq1 \mgmtsoc_load_storage_reg[10]  ( .D(n3424), .CP(n6084), .Q(
        csrbank10_load0_w[10]) );
  dfnrq1 \mgmtsoc_value_reg[10]  ( .D(N5410), .CP(n6102), .Q(mgmtsoc_value[10]) );
  dfnrq1 \mgmtsoc_value_status_reg[10]  ( .D(n3490), .CP(n6124), .Q(
        csrbank10_value_w[10]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[10]  ( .D(N4704), .CP(n6092), .Q(
        interface10_bank_bus_dat_r[10]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[10]  ( .D(n3317), .CP(n6093), .Q(
        csrbank0_scratch0_w[10]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[10]  ( .D(N4109), .CP(n6095), .Q(
        interface0_bank_bus_dat_r[10]) );
  dfnrq1 \memdat_3_reg[3]  ( .D(n3738), .CP(n6095), .Q(
        uart_rx_fifo_fifo_out_payload_data[3]) );
  dfnrq1 \interface11_bank_bus_dat_r_reg[3]  ( .D(N4775), .CP(n6102), .Q(
        interface11_bank_bus_dat_r[3]) );
  dfnrq1 \dbg_uart_data_reg[3]  ( .D(n3280), .CP(n6084), .Q(
        dbg_uart_wishbone_dat_w[3]) );
  dfnrq1 \spi_master_mosi_storage_reg[3]  ( .D(n4542), .CP(n6124), .Q(
        spi_master_mosi[3]) );
  dfnrq1 \spi_master_mosi_data_reg[3]  ( .D(n3690), .CP(n6092), .Q(
        spi_master_mosi_data[3]) );
  dfnrq1 \la_out_storage_reg[3]  ( .D(n4477), .CP(n6093), .Q(n131) );
  dfnrq1 \la_out_storage_reg[35]  ( .D(n4445), .CP(n6096), .Q(n99) );
  dfnrq1 \la_out_storage_reg[67]  ( .D(n4413), .CP(n6095), .Q(n67) );
  dfnrq1 \la_out_storage_reg[99]  ( .D(n4381), .CP(n6092), .Q(n35) );
  dfnrq1 \la_oe_storage_reg[3]  ( .D(n4349), .CP(n6092), .Q(csrbank6_oe0_w[3])
         );
  dfnrq1 \la_oe_storage_reg[35]  ( .D(n4317), .CP(n6092), .Q(csrbank6_oe1_w[3]) );
  dfnrq1 \la_oe_storage_reg[67]  ( .D(n4285), .CP(n6092), .Q(csrbank6_oe2_w[3]) );
  dfnrq1 \la_oe_storage_reg[99]  ( .D(n4253), .CP(n6092), .Q(csrbank6_oe3_w[3]) );
  dfnrq1 \la_ien_storage_reg[3]  ( .D(n4221), .CP(n6092), .Q(
        csrbank6_ien0_w[3]) );
  dfnrq1 \la_ien_storage_reg[35]  ( .D(n4189), .CP(n6092), .Q(
        csrbank6_ien1_w[3]) );
  dfnrq1 \la_ien_storage_reg[67]  ( .D(n4157), .CP(n6092), .Q(
        csrbank6_ien2_w[3]) );
  dfnrq1 \la_ien_storage_reg[99]  ( .D(n4125), .CP(n6093), .Q(
        csrbank6_ien3_w[3]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[3]  ( .D(N4466), .CP(n6093), .Q(
        interface6_bank_bus_dat_r[3]) );
  dfnrq1 \storage_reg[15][3]  ( .D(n4036), .CP(n6093), .Q(\storage[15][3] ) );
  dfnrq1 \storage_reg[14][3]  ( .D(n4028), .CP(n6093), .Q(\storage[14][3] ) );
  dfnrq1 \storage_reg[13][3]  ( .D(n4020), .CP(n6093), .Q(\storage[13][3] ) );
  dfnrq1 \storage_reg[12][3]  ( .D(n4012), .CP(n6093), .Q(\storage[12][3] ) );
  dfnrq1 \storage_reg[11][3]  ( .D(n4004), .CP(n6093), .Q(\storage[11][3] ) );
  dfnrq1 \storage_reg[10][3]  ( .D(n3996), .CP(n6093), .Q(\storage[10][3] ) );
  dfnrq1 \storage_reg[9][3]  ( .D(n3988), .CP(n6074), .Q(\storage[9][3] ) );
  dfnrq1 \storage_reg[8][3]  ( .D(n3980), .CP(n6099), .Q(\storage[8][3] ) );
  dfnrq1 \storage_reg[7][3]  ( .D(n3972), .CP(n6074), .Q(\storage[7][3] ) );
  dfnrq1 \storage_reg[6][3]  ( .D(n3964), .CP(n6099), .Q(\storage[6][3] ) );
  dfnrq1 \storage_reg[5][3]  ( .D(n3956), .CP(n6074), .Q(\storage[5][3] ) );
  dfnrq1 \storage_reg[4][3]  ( .D(n3948), .CP(n6074), .Q(\storage[4][3] ) );
  dfnrq1 \storage_reg[3][3]  ( .D(n3940), .CP(n6074), .Q(\storage[3][3] ) );
  dfnrq1 \storage_reg[2][3]  ( .D(n3932), .CP(n6074), .Q(\storage[2][3] ) );
  dfnrq1 \storage_reg[1][3]  ( .D(n3924), .CP(n6088), .Q(\storage[1][3] ) );
  dfnrq1 \storage_reg[0][3]  ( .D(n3916), .CP(n6089), .Q(\storage[0][3] ) );
  dfnrq1 \memdat_1_reg[3]  ( .D(n3894), .CP(n6024), .Q(
        uart_tx_fifo_fifo_out_payload_data[3]) );
  dfnrq1 \spimaster_storage_reg[3]  ( .D(n3717), .CP(n6101), .Q(
        spi_master_clk_divider0[3]) );
  dfnrq1 \spi_master_cs_storage_reg[3]  ( .D(n3678), .CP(n6045), .Q(
        csrbank9_cs0_w[3]) );
  dfnrq1 \spi_master_control_storage_reg[3]  ( .D(n3659), .CP(n6044), .Q(
        csrbank9_control0_w[3]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[3]  ( .D(N4588), .CP(n6039), .Q(
        interface9_bank_bus_dat_r[3]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[3]  ( .D(n3599), .CP(
        n6107), .Q(mgmtsoc_port_master_user_port_sink_payload_data[3]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[3]  ( .D(n3556), .CP(n6107), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_len[3]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_len_reg[3]  ( .D(n3567), .CP(
        n6108), .Q(mgmtsoc_port_master_user_port_sink_payload_len[3]) );
  dfnrq1 \mgmtsoc_litespimmap_storage_reg[3]  ( .D(n3531), .CP(n6107), .Q(
        mgmtsoc_litespimmap_spi_dummy_bits[3]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[3]  ( .D(N4246), .CP(n6107), .Q(
        interface3_bank_bus_dat_r[3]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_storage_reg[3]  ( .D(n3508), .CP(n6107), 
        .Q(mgmtsoc_litespisdrphycore_div[3]) );
  dfnrq1 \interface4_bank_bus_dat_r_reg[3]  ( .D(N4295), .CP(n6107), .Q(
        interface4_bank_bus_dat_r[3]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[3]  ( .D(n3463), .CP(n6107), .Q(
        csrbank10_reload0_w[3]) );
  dfnrq1 \mgmtsoc_load_storage_reg[3]  ( .D(n3431), .CP(n6107), .Q(
        csrbank10_load0_w[3]) );
  dfnrq1 \mgmtsoc_value_reg[3]  ( .D(N5403), .CP(n6107), .Q(mgmtsoc_value[3])
         );
  dfnrq1 \mgmtsoc_value_status_reg[3]  ( .D(n3497), .CP(n6107), .Q(
        csrbank10_value_w[3]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[3]  ( .D(N4697), .CP(n6062), .Q(
        interface10_bank_bus_dat_r[3]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[3]  ( .D(n3324), .CP(n6108), .Q(
        csrbank0_scratch0_w[3]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[3]  ( .D(N4102), .CP(n6129), .Q(
        interface0_bank_bus_dat_r[3]) );
  dfnrq1 \memdat_3_reg[4]  ( .D(n3736), .CP(n6106), .Q(
        uart_rx_fifo_fifo_out_payload_data[4]) );
  dfnrq1 \interface11_bank_bus_dat_r_reg[4]  ( .D(N4776), .CP(n6105), .Q(
        interface11_bank_bus_dat_r[4]) );
  dfnrq1 \memdat_3_reg[5]  ( .D(n3734), .CP(n6129), .Q(
        uart_rx_fifo_fifo_out_payload_data[5]) );
  dfnrq1 \interface11_bank_bus_dat_r_reg[5]  ( .D(N4777), .CP(n6063), .Q(
        interface11_bank_bus_dat_r[5]) );
  dfnrq1 \dbg_uart_data_reg[5]  ( .D(n3278), .CP(n6129), .Q(
        dbg_uart_wishbone_dat_w[5]) );
  dfnrq1 \spi_master_mosi_storage_reg[5]  ( .D(n4540), .CP(n6108), .Q(
        spi_master_mosi[5]) );
  dfnrq1 \spi_master_mosi_data_reg[5]  ( .D(n3688), .CP(n6108), .Q(
        spi_master_mosi_data[5]) );
  dfnrq1 \la_out_storage_reg[5]  ( .D(n4475), .CP(n6108), .Q(n129) );
  dfnrq1 \la_out_storage_reg[37]  ( .D(n4443), .CP(n6108), .Q(n97) );
  dfnrq1 \la_out_storage_reg[69]  ( .D(n4411), .CP(n6108), .Q(n65) );
  dfnrq1 \la_out_storage_reg[101]  ( .D(n4379), .CP(n6108), .Q(n33) );
  dfnrq1 \la_oe_storage_reg[5]  ( .D(n4347), .CP(n6108), .Q(csrbank6_oe0_w[5])
         );
  dfnrq1 \la_oe_storage_reg[37]  ( .D(n4315), .CP(n6108), .Q(csrbank6_oe1_w[5]) );
  dfnrq1 \la_oe_storage_reg[69]  ( .D(n4283), .CP(n6081), .Q(csrbank6_oe2_w[5]) );
  dfnrq1 \la_oe_storage_reg[101]  ( .D(n4251), .CP(n6097), .Q(
        csrbank6_oe3_w[5]) );
  dfnrq1 \la_ien_storage_reg[5]  ( .D(n4219), .CP(n6076), .Q(
        csrbank6_ien0_w[5]) );
  dfnrq1 \la_ien_storage_reg[37]  ( .D(n4187), .CP(n6089), .Q(
        csrbank6_ien1_w[5]) );
  dfnrq1 \la_ien_storage_reg[69]  ( .D(n4155), .CP(n6040), .Q(
        csrbank6_ien2_w[5]) );
  dfnrq1 \la_ien_storage_reg[101]  ( .D(n4123), .CP(n6087), .Q(
        csrbank6_ien3_w[5]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[5]  ( .D(N4468), .CP(n6079), .Q(
        interface6_bank_bus_dat_r[5]) );
  dfnrq1 \storage_reg[15][5]  ( .D(n4034), .CP(n6033), .Q(\storage[15][5] ) );
  dfnrq1 \storage_reg[14][5]  ( .D(n4026), .CP(n6109), .Q(\storage[14][5] ) );
  dfnrq1 \storage_reg[13][5]  ( .D(n4018), .CP(n6129), .Q(\storage[13][5] ) );
  dfnrq1 \storage_reg[12][5]  ( .D(n4010), .CP(n6110), .Q(\storage[12][5] ) );
  dfnrq1 \storage_reg[11][5]  ( .D(n4002), .CP(n6096), .Q(\storage[11][5] ) );
  dfnrq1 \storage_reg[10][5]  ( .D(n3994), .CP(n6024), .Q(\storage[10][5] ) );
  dfnrq1 \storage_reg[9][5]  ( .D(n3986), .CP(n6109), .Q(\storage[9][5] ) );
  dfnrq1 \storage_reg[8][5]  ( .D(n3978), .CP(n6103), .Q(\storage[8][5] ) );
  dfnrq1 \storage_reg[7][5]  ( .D(n3970), .CP(n6129), .Q(\storage[7][5] ) );
  dfnrq1 \storage_reg[6][5]  ( .D(n3962), .CP(n6109), .Q(\storage[6][5] ) );
  dfnrq1 \storage_reg[5][5]  ( .D(n3954), .CP(n6109), .Q(\storage[5][5] ) );
  dfnrq1 \storage_reg[4][5]  ( .D(n3946), .CP(n6109), .Q(\storage[4][5] ) );
  dfnrq1 \storage_reg[3][5]  ( .D(n3938), .CP(n6109), .Q(\storage[3][5] ) );
  dfnrq1 \storage_reg[2][5]  ( .D(n3930), .CP(n6109), .Q(\storage[2][5] ) );
  dfnrq1 \storage_reg[1][5]  ( .D(n3922), .CP(n6109), .Q(\storage[1][5] ) );
  dfnrq1 \storage_reg[0][5]  ( .D(n3914), .CP(n6109), .Q(\storage[0][5] ) );
  dfnrq1 \memdat_1_reg[5]  ( .D(n3896), .CP(n6109), .Q(
        uart_tx_fifo_fifo_out_payload_data[5]) );
  dfnrq1 \uart_phy_tx_data_reg[5]  ( .D(n3886), .CP(n6067), .Q(
        uart_phy_tx_data[5]) );
  dfnrq1 \spimaster_storage_reg[5]  ( .D(n3715), .CP(n6110), .Q(
        spi_master_clk_divider0[5]) );
  dfnrq1 \spi_master_cs_storage_reg[5]  ( .D(n3676), .CP(n6060), .Q(
        csrbank9_cs0_w[5]) );
  dfnrq1 \spi_master_control_storage_reg[5]  ( .D(n3657), .CP(n6107), .Q(
        csrbank9_control0_w[5]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[5]  ( .D(N4590), .CP(n6103), .Q(
        interface9_bank_bus_dat_r[5]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[5]  ( .D(n3597), .CP(
        n6129), .Q(mgmtsoc_port_master_user_port_sink_payload_data[5]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[5]  ( .D(n3554), .CP(n6110), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_len[5]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_len_reg[5]  ( .D(n3565), .CP(
        n6101), .Q(mgmtsoc_port_master_user_port_sink_payload_len[5]) );
  dfnrq1 \mgmtsoc_litespimmap_storage_reg[5]  ( .D(n3529), .CP(n6108), .Q(
        mgmtsoc_litespimmap_spi_dummy_bits[5]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[5]  ( .D(N4248), .CP(n6029), .Q(
        interface3_bank_bus_dat_r[5]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_storage_reg[5]  ( .D(n3506), .CP(n6129), 
        .Q(mgmtsoc_litespisdrphycore_div[5]) );
  dfnrq1 \interface4_bank_bus_dat_r_reg[5]  ( .D(N4297), .CP(n6095), .Q(
        interface4_bank_bus_dat_r[5]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[5]  ( .D(n3461), .CP(n6129), .Q(
        csrbank10_reload0_w[5]) );
  dfnrq1 \mgmtsoc_load_storage_reg[5]  ( .D(n3429), .CP(n6129), .Q(
        csrbank10_load0_w[5]) );
  dfnrq1 \mgmtsoc_value_reg[5]  ( .D(N5405), .CP(n6104), .Q(mgmtsoc_value[5])
         );
  dfnrq1 \mgmtsoc_value_status_reg[5]  ( .D(n3495), .CP(n6110), .Q(
        csrbank10_value_w[5]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[5]  ( .D(N4699), .CP(n6110), .Q(
        interface10_bank_bus_dat_r[5]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[5]  ( .D(n3322), .CP(n6110), .Q(
        csrbank0_scratch0_w[5]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[5]  ( .D(N4104), .CP(n6110), .Q(
        interface0_bank_bus_dat_r[5]) );
  dfnrq1 \memdat_3_reg[6]  ( .D(n3732), .CP(n6110), .Q(
        uart_rx_fifo_fifo_out_payload_data[6]) );
  dfnrq1 \interface11_bank_bus_dat_r_reg[6]  ( .D(N4778), .CP(n6110), .Q(
        interface11_bank_bus_dat_r[6]) );
  dfnrq1 \memdat_3_reg[7]  ( .D(n3730), .CP(n6110), .Q(
        uart_rx_fifo_fifo_out_payload_data[7]) );
  dfnrq1 \interface11_bank_bus_dat_r_reg[7]  ( .D(N4779), .CP(n6110), .Q(
        interface11_bank_bus_dat_r[7]) );
  dfnrq1 \mgmtsoc_reset_storage_reg[1]  ( .D(n3294), .CP(n6056), .Q(
        csrbank0_reset0_w[1]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[1]  ( .D(N4100), .CP(n6091), .Q(
        interface0_bank_bus_dat_r[1]) );
  dfnrq1 \dbg_uart_data_reg[9]  ( .D(n3274), .CP(n6090), .Q(
        dbg_uart_wishbone_dat_w[9]) );
  dfnrq1 \la_out_storage_reg[9]  ( .D(n4471), .CP(n6094), .Q(n125) );
  dfnrq1 \la_out_storage_reg[41]  ( .D(n4439), .CP(n6048), .Q(n93) );
  dfnrq1 \la_out_storage_reg[73]  ( .D(n4407), .CP(n6041), .Q(n61) );
  dfnrq1 \la_out_storage_reg[105]  ( .D(n4375), .CP(n6092), .Q(n29) );
  dfnrq1 \la_oe_storage_reg[9]  ( .D(n4343), .CP(n6093), .Q(csrbank6_oe0_w[9])
         );
  dfnrq1 \la_oe_storage_reg[41]  ( .D(n4311), .CP(n6110), .Q(csrbank6_oe1_w[9]) );
  dfnrq1 \la_oe_storage_reg[73]  ( .D(n4279), .CP(n6109), .Q(csrbank6_oe2_w[9]) );
  dfnrq1 \la_oe_storage_reg[105]  ( .D(n4247), .CP(n6107), .Q(
        csrbank6_oe3_w[9]) );
  dfnrq1 \la_ien_storage_reg[9]  ( .D(n4215), .CP(n6106), .Q(
        csrbank6_ien0_w[9]) );
  dfnrq1 \la_ien_storage_reg[41]  ( .D(n4183), .CP(n6105), .Q(
        csrbank6_ien1_w[9]) );
  dfnrq1 \la_ien_storage_reg[73]  ( .D(n4151), .CP(n6104), .Q(
        csrbank6_ien2_w[9]) );
  dfnrq1 \la_ien_storage_reg[105]  ( .D(n4119), .CP(n6103), .Q(
        csrbank6_ien3_w[9]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[9]  ( .D(N4472), .CP(n6129), .Q(
        interface6_bank_bus_dat_r[9]) );
  dfnrq1 \spimaster_storage_reg[9]  ( .D(n3711), .CP(n6069), .Q(
        spi_master_clk_divider0[9]) );
  dfnrq1 \spi_master_cs_storage_reg[9]  ( .D(n3672), .CP(n6129), .Q(
        csrbank9_cs0_w[9]) );
  dfnrq1 \spi_master_control_storage_reg[9]  ( .D(n3653), .CP(n6068), .Q(
        spi_master_length0[1]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[9]  ( .D(N4594), .CP(n6129), .Q(
        interface9_bank_bus_dat_r[9]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[9]  ( .D(n3593), .CP(
        n6066), .Q(mgmtsoc_port_master_user_port_sink_payload_data[9]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[9]  ( .D(n3550), .CP(n6109), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_width[1]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[9]  ( .D(N4252), .CP(n6073), .Q(
        interface3_bank_bus_dat_r[9]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_width_reg[1]  ( .D(n3563), 
        .CP(n6110), .Q(mgmtsoc_port_master_user_port_sink_payload_width[1]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[9]  ( .D(n3457), .CP(n6072), .Q(
        csrbank10_reload0_w[9]) );
  dfnrq1 \mgmtsoc_load_storage_reg[9]  ( .D(n3425), .CP(n6106), .Q(
        csrbank10_load0_w[9]) );
  dfnrq1 \mgmtsoc_value_reg[9]  ( .D(N5409), .CP(n6071), .Q(mgmtsoc_value[9])
         );
  dfnrq1 \mgmtsoc_value_status_reg[9]  ( .D(n3491), .CP(n6108), .Q(
        csrbank10_value_w[9]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[9]  ( .D(N4703), .CP(n6070), .Q(
        interface10_bank_bus_dat_r[9]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[9]  ( .D(n3318), .CP(n6107), .Q(
        csrbank0_scratch0_w[9]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[9]  ( .D(N4108), .CP(n6064), .Q(
        interface0_bank_bus_dat_r[9]) );
  dfnrq1 \spi_master_miso_reg[0]  ( .D(n3646), .CP(n6103), .Q(
        spi_master_miso_status[0]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[0]  ( .D(N4585), .CP(n6065), .Q(
        interface9_bank_bus_dat_r[0]) );
  dfnrq1 \la_out_storage_reg[4]  ( .D(n4476), .CP(n6104), .Q(n130) );
  dfnrq1 \la_out_storage_reg[36]  ( .D(n4444), .CP(n6108), .Q(n98) );
  dfnrq1 \la_out_storage_reg[68]  ( .D(n4412), .CP(n6129), .Q(n66) );
  dfnrq1 \la_out_storage_reg[100]  ( .D(n4380), .CP(n6109), .Q(n34) );
  dfnrq1 \la_oe_storage_reg[4]  ( .D(n4348), .CP(n6122), .Q(csrbank6_oe0_w[4])
         );
  dfnrq1 \la_oe_storage_reg[36]  ( .D(n4316), .CP(n6112), .Q(csrbank6_oe1_w[4]) );
  dfnrq1 \la_oe_storage_reg[68]  ( .D(n4284), .CP(n6088), .Q(csrbank6_oe2_w[4]) );
  dfnrq1 \la_oe_storage_reg[100]  ( .D(n4252), .CP(n6059), .Q(
        csrbank6_oe3_w[4]) );
  dfnrq1 \la_ien_storage_reg[4]  ( .D(n4220), .CP(n6110), .Q(
        csrbank6_ien0_w[4]) );
  dfnrq1 \la_ien_storage_reg[36]  ( .D(n4188), .CP(n6102), .Q(
        csrbank6_ien1_w[4]) );
  dfnrq1 \la_ien_storage_reg[68]  ( .D(n4156), .CP(n6084), .Q(
        csrbank6_ien2_w[4]) );
  dfnrq1 \la_ien_storage_reg[100]  ( .D(n4124), .CP(n6104), .Q(
        csrbank6_ien3_w[4]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[4]  ( .D(N4467), .CP(n6098), .Q(
        interface6_bank_bus_dat_r[4]) );
  dfnrq1 \storage_reg[15][4]  ( .D(n4035), .CP(n6098), .Q(\storage[15][4] ) );
  dfnrq1 \storage_reg[14][4]  ( .D(n4027), .CP(n6099), .Q(\storage[14][4] ) );
  dfnrq1 \storage_reg[13][4]  ( .D(n4019), .CP(n6099), .Q(\storage[13][4] ) );
  dfnrq1 \storage_reg[12][4]  ( .D(n4011), .CP(n6099), .Q(\storage[12][4] ) );
  dfnrq1 \storage_reg[11][4]  ( .D(n4003), .CP(n6099), .Q(\storage[11][4] ) );
  dfnrq1 \storage_reg[10][4]  ( .D(n3995), .CP(n6099), .Q(\storage[10][4] ) );
  dfnrq1 \storage_reg[9][4]  ( .D(n3987), .CP(n6099), .Q(\storage[9][4] ) );
  dfnrq1 \storage_reg[8][4]  ( .D(n3979), .CP(n6099), .Q(\storage[8][4] ) );
  dfnrq1 \storage_reg[7][4]  ( .D(n3971), .CP(n6099), .Q(\storage[7][4] ) );
  dfnrq1 \storage_reg[6][4]  ( .D(n3963), .CP(n6100), .Q(\storage[6][4] ) );
  dfnrq1 \storage_reg[5][4]  ( .D(n3955), .CP(n6100), .Q(\storage[5][4] ) );
  dfnrq1 \storage_reg[4][4]  ( .D(n3947), .CP(n6100), .Q(\storage[4][4] ) );
  dfnrq1 \storage_reg[3][4]  ( .D(n3939), .CP(n6100), .Q(\storage[3][4] ) );
  dfnrq1 \storage_reg[2][4]  ( .D(n3931), .CP(n6100), .Q(\storage[2][4] ) );
  dfnrq1 \storage_reg[1][4]  ( .D(n3923), .CP(n6100), .Q(\storage[1][4] ) );
  dfnrq1 \storage_reg[0][4]  ( .D(n3915), .CP(n6100), .Q(\storage[0][4] ) );
  dfnrq1 \memdat_1_reg[4]  ( .D(n3895), .CP(n6100), .Q(
        uart_tx_fifo_fifo_out_payload_data[4]) );
  dfnrq1 \uart_phy_tx_data_reg[4]  ( .D(n3887), .CP(n6086), .Q(
        uart_phy_tx_data[4]) );
  dfnrq1 \uart_phy_tx_data_reg[3]  ( .D(n3888), .CP(n6024), .Q(
        uart_phy_tx_data[3]) );
  dfnrq1 \uart_phy_tx_data_reg[2]  ( .D(n3889), .CP(n6125), .Q(
        uart_phy_tx_data[2]) );
  dfnrq1 \uart_phy_tx_data_reg[1]  ( .D(n3890), .CP(n6093), .Q(
        uart_phy_tx_data[1]) );
  dfnrq1 \uart_phy_tx_data_reg[0]  ( .D(n3891), .CP(n6124), .Q(
        uart_phy_tx_data[0]) );
  dfnrq1 sys_uart_tx_reg ( .D(n3883), .CP(n6103), .Q(sys_uart_tx) );
  dfnrq1 \spimaster_storage_reg[4]  ( .D(n3716), .CP(n6110), .Q(
        spi_master_clk_divider0[4]) );
  dfnrq1 \spi_master_cs_storage_reg[4]  ( .D(n3677), .CP(n6107), .Q(
        csrbank9_cs0_w[4]) );
  dfnrq1 \spi_master_control_storage_reg[4]  ( .D(n3658), .CP(n6101), .Q(
        csrbank9_control0_w[4]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[4]  ( .D(N4589), .CP(n6101), .Q(
        interface9_bank_bus_dat_r[4]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[4]  ( .D(n3598), .CP(
        n6101), .Q(mgmtsoc_port_master_user_port_sink_payload_data[4]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[4]  ( .D(n3555), .CP(n6101), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_len[4]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_len_reg[4]  ( .D(n3566), .CP(
        n6101), .Q(mgmtsoc_port_master_user_port_sink_payload_len[4]) );
  dfnrq1 \mgmtsoc_litespimmap_storage_reg[4]  ( .D(n3530), .CP(n6101), .Q(
        mgmtsoc_litespimmap_spi_dummy_bits[4]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[4]  ( .D(N4247), .CP(n6101), .Q(
        interface3_bank_bus_dat_r[4]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_storage_reg[4]  ( .D(n3507), .CP(n6101), 
        .Q(mgmtsoc_litespisdrphycore_div[4]) );
  dfnrq1 \interface4_bank_bus_dat_r_reg[4]  ( .D(N4296), .CP(n6102), .Q(
        interface4_bank_bus_dat_r[4]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[4]  ( .D(n3462), .CP(n6102), .Q(
        csrbank10_reload0_w[4]) );
  dfnrq1 \mgmtsoc_load_storage_reg[4]  ( .D(n3430), .CP(n6102), .Q(
        csrbank10_load0_w[4]) );
  dfnrq1 \mgmtsoc_value_reg[4]  ( .D(N5404), .CP(n6102), .Q(mgmtsoc_value[4])
         );
  dfnrq1 \mgmtsoc_value_status_reg[4]  ( .D(n3496), .CP(n6102), .Q(
        csrbank10_value_w[4]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[4]  ( .D(N4698), .CP(n6102), .Q(
        interface10_bank_bus_dat_r[4]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[4]  ( .D(n3323), .CP(n6102), .Q(
        csrbank0_scratch0_w[4]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[4]  ( .D(N4103), .CP(n6102), .Q(
        interface0_bank_bus_dat_r[4]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_mask_reg[0]  ( .D(n3560), .CP(
        n6090), .Q(\mgmtsoc_port_master_user_port_sink_payload_mask[0] ) );
  dfnrq1 flash_io0_oeb_reg ( .D(n4547), .CP(n6104), .Q(flash_io0_oeb) );
  dfnrq1 \mgmtsoc_reload_storage_reg[6]  ( .D(n3460), .CP(n6084), .Q(
        csrbank10_reload0_w[6]) );
  dfnrq1 \mgmtsoc_load_storage_reg[6]  ( .D(n3428), .CP(n6124), .Q(
        csrbank10_load0_w[6]) );
  dfnrq1 \mgmtsoc_value_reg[6]  ( .D(N5406), .CP(n6107), .Q(mgmtsoc_value[6])
         );
  dfnrq1 \mgmtsoc_value_status_reg[6]  ( .D(n3494), .CP(n6057), .Q(
        csrbank10_value_w[6]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[6]  ( .D(N4700), .CP(n6125), .Q(
        interface10_bank_bus_dat_r[6]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[6]  ( .D(n3321), .CP(n6086), .Q(
        csrbank0_scratch0_w[6]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[6]  ( .D(N4105), .CP(n6103), .Q(
        interface0_bank_bus_dat_r[6]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_cnt_reg[1]  ( .D(n3127), .CP(n6103), 
        .Q(mgmtsoc_litespisdrphycore_sr_cnt[1]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_cnt_reg[0]  ( .D(n3126), .CP(n6103), 
        .Q(mgmtsoc_litespisdrphycore_sr_cnt[0]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_cnt_reg[2]  ( .D(n3125), .CP(n6103), 
        .Q(mgmtsoc_litespisdrphycore_sr_cnt[2]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_cnt_reg[3]  ( .D(n3124), .CP(n6103), 
        .Q(mgmtsoc_litespisdrphycore_sr_cnt[3]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_cnt_reg[4]  ( .D(n3123), .CP(n6103), 
        .Q(mgmtsoc_litespisdrphycore_sr_cnt[4]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_cnt_reg[5]  ( .D(n3122), .CP(n6103), 
        .Q(mgmtsoc_litespisdrphycore_sr_cnt[5]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_cnt_reg[6]  ( .D(n3121), .CP(n6103), 
        .Q(mgmtsoc_litespisdrphycore_sr_cnt[6]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[7]  ( .D(n3459), .CP(n6104), .Q(
        csrbank10_reload0_w[7]) );
  dfnrq1 \mgmtsoc_load_storage_reg[7]  ( .D(n3427), .CP(n6104), .Q(
        csrbank10_load0_w[7]) );
  dfnrq1 \mgmtsoc_value_reg[7]  ( .D(N5407), .CP(n6104), .Q(mgmtsoc_value[7])
         );
  dfnrq1 \mgmtsoc_value_status_reg[7]  ( .D(n3493), .CP(n6104), .Q(
        csrbank10_value_w[7]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[7]  ( .D(N4701), .CP(n6104), .Q(
        interface10_bank_bus_dat_r[7]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[7]  ( .D(n3320), .CP(n6104), .Q(
        csrbank0_scratch0_w[7]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[7]  ( .D(N4106), .CP(n6104), .Q(
        interface0_bank_bus_dat_r[7]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[0]  ( .D(n3159), .CP(n6105), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[0]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[1]  ( .D(n3128), .CP(n6105), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[1]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[2]  ( .D(n3129), .CP(n6105), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[2]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[3]  ( .D(n3130), .CP(n6105), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[3]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[4]  ( .D(n3131), .CP(n6105), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[4]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[5]  ( .D(n3132), .CP(n6105), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[5]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[6]  ( .D(n3133), .CP(n6105), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[6]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[7]  ( .D(n3134), .CP(n6105), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[7]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[8]  ( .D(n3135), .CP(n6106), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[8]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[9]  ( .D(n3136), .CP(n6106), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[9]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[10]  ( .D(n3137), .CP(n6106), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[10]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[11]  ( .D(n3138), .CP(n6106), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[11]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[11]  ( .D(n3455), .CP(n6106), .Q(
        csrbank10_reload0_w[11]) );
  dfnrq1 \mgmtsoc_load_storage_reg[11]  ( .D(n3423), .CP(n6106), .Q(
        csrbank10_load0_w[11]) );
  dfnrq1 \mgmtsoc_value_reg[11]  ( .D(N5411), .CP(n6106), .Q(mgmtsoc_value[11]) );
  dfnrq1 \mgmtsoc_value_status_reg[11]  ( .D(n3489), .CP(n6106), .Q(
        csrbank10_value_w[11]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[11]  ( .D(N4705), .CP(n6110), .Q(
        interface10_bank_bus_dat_r[11]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[11]  ( .D(n3316), .CP(n6086), .Q(
        csrbank0_scratch0_w[11]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[11]  ( .D(N4110), .CP(n6119), .Q(
        interface0_bank_bus_dat_r[11]) );
  dfnrq1 \dbg_uart_data_reg[12]  ( .D(n3271), .CP(n6109), .Q(
        dbg_uart_wishbone_dat_w[12]) );
  dfnrq1 \la_out_storage_reg[12]  ( .D(n4468), .CP(n6129), .Q(n122) );
  dfnrq1 \la_out_storage_reg[44]  ( .D(n4436), .CP(n6106), .Q(n90) );
  dfnrq1 \la_out_storage_reg[76]  ( .D(n4404), .CP(n6105), .Q(n58) );
  dfnrq1 \la_out_storage_reg[108]  ( .D(n4372), .CP(n6108), .Q(n26) );
  dfnrq1 \la_oe_storage_reg[12]  ( .D(n4340), .CP(n6110), .Q(
        csrbank6_oe0_w[12]) );
  dfnrq1 \la_oe_storage_reg[44]  ( .D(n4308), .CP(n6108), .Q(
        csrbank6_oe1_w[12]) );
  dfnrq1 \la_oe_storage_reg[76]  ( .D(n4276), .CP(n6085), .Q(
        csrbank6_oe2_w[12]) );
  dfnrq1 \la_oe_storage_reg[108]  ( .D(n4244), .CP(n6108), .Q(
        csrbank6_oe3_w[12]) );
  dfnrq1 \la_ien_storage_reg[12]  ( .D(n4212), .CP(n6103), .Q(
        csrbank6_ien0_w[12]) );
  dfnrq1 \la_ien_storage_reg[44]  ( .D(n4180), .CP(n6108), .Q(
        csrbank6_ien1_w[12]) );
  dfnrq1 \la_ien_storage_reg[76]  ( .D(n4148), .CP(n6104), .Q(
        csrbank6_ien2_w[12]) );
  dfnrq1 \la_ien_storage_reg[108]  ( .D(n4116), .CP(n6108), .Q(
        csrbank6_ien3_w[12]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[12]  ( .D(N4475), .CP(n6107), .Q(
        interface6_bank_bus_dat_r[12]) );
  dfnrq1 \spimaster_storage_reg[12]  ( .D(n3708), .CP(n6104), .Q(
        spi_master_clk_divider0[12]) );
  dfnrq1 \spi_master_cs_storage_reg[12]  ( .D(n3669), .CP(n6103), .Q(
        csrbank9_cs0_w[12]) );
  dfnrq1 \spi_master_control_storage_reg[12]  ( .D(n3650), .CP(n6109), .Q(
        spi_master_length0[4]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[12]  ( .D(N4597), .CP(n6106), .Q(
        interface9_bank_bus_dat_r[12]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[12]  ( .D(n3590), 
        .CP(n6025), .Q(mgmtsoc_port_master_user_port_sink_payload_data[12]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[12]  ( .D(n3139), .CP(n6106), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[12]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[12]  ( .D(n3547), .CP(n6107), 
        .Q(csrbank3_master_phyconfig0_w[12]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[12]  ( .D(N4255), .CP(n6106), .Q(
        interface3_bank_bus_dat_r[12]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[12]  ( .D(n3454), .CP(n6026), .Q(
        csrbank10_reload0_w[12]) );
  dfnrq1 \mgmtsoc_load_storage_reg[12]  ( .D(n3422), .CP(n6107), .Q(
        csrbank10_load0_w[12]) );
  dfnrq1 \mgmtsoc_value_reg[12]  ( .D(N5412), .CP(n6104), .Q(mgmtsoc_value[12]) );
  dfnrq1 \mgmtsoc_value_status_reg[12]  ( .D(n3488), .CP(n6108), .Q(
        csrbank10_value_w[12]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[12]  ( .D(N4706), .CP(n6109), .Q(
        interface10_bank_bus_dat_r[12]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[12]  ( .D(n3315), .CP(n6129), .Q(
        csrbank0_scratch0_w[12]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[12]  ( .D(N4111), .CP(n6106), .Q(
        interface0_bank_bus_dat_r[12]) );
  dfnrq1 \dbg_uart_data_reg[13]  ( .D(n3270), .CP(n6103), .Q(
        dbg_uart_wishbone_dat_w[13]) );
  dfnrq1 \la_out_storage_reg[13]  ( .D(n4467), .CP(n6129), .Q(n121) );
  dfnrq1 \la_out_storage_reg[45]  ( .D(n4435), .CP(n6057), .Q(n89) );
  dfnrq1 \la_out_storage_reg[77]  ( .D(n4403), .CP(n6104), .Q(n57) );
  dfnrq1 \la_out_storage_reg[109]  ( .D(n4371), .CP(n6104), .Q(n25) );
  dfnrq1 \la_oe_storage_reg[13]  ( .D(n4339), .CP(n6103), .Q(
        csrbank6_oe0_w[13]) );
  dfnrq1 \la_oe_storage_reg[45]  ( .D(n4307), .CP(n6078), .Q(
        csrbank6_oe1_w[13]) );
  dfnrq1 \la_oe_storage_reg[77]  ( .D(n4275), .CP(n6069), .Q(
        csrbank6_oe2_w[13]) );
  dfnrq1 \la_oe_storage_reg[109]  ( .D(n4243), .CP(n6117), .Q(
        csrbank6_oe3_w[13]) );
  dfnrq1 \la_ien_storage_reg[13]  ( .D(n4211), .CP(n6068), .Q(
        csrbank6_ien0_w[13]) );
  dfnrq1 \la_ien_storage_reg[45]  ( .D(n4179), .CP(n6066), .Q(
        csrbank6_ien1_w[13]) );
  dfnrq1 \la_ien_storage_reg[77]  ( .D(n4147), .CP(n6117), .Q(
        csrbank6_ien2_w[13]) );
  dfnrq1 \la_ien_storage_reg[109]  ( .D(n4115), .CP(n6068), .Q(
        csrbank6_ien3_w[13]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[13]  ( .D(N4476), .CP(n6067), .Q(
        interface6_bank_bus_dat_r[13]) );
  dfnrq1 \spimaster_storage_reg[13]  ( .D(n3707), .CP(n6070), .Q(
        spi_master_clk_divider0[13]) );
  dfnrq1 \spi_master_cs_storage_reg[13]  ( .D(n3668), .CP(n6070), .Q(
        csrbank9_cs0_w[13]) );
  dfnrq1 \spi_master_control_storage_reg[13]  ( .D(n3649), .CP(n6070), .Q(
        spi_master_length0[5]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[13]  ( .D(N4598), .CP(n6070), .Q(
        interface9_bank_bus_dat_r[13]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[13]  ( .D(n3589), 
        .CP(n6070), .Q(mgmtsoc_port_master_user_port_sink_payload_data[13]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[13]  ( .D(n3140), .CP(n6070), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[13]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[13]  ( .D(n3546), .CP(n6070), 
        .Q(csrbank3_master_phyconfig0_w[13]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[13]  ( .D(N4256), .CP(n6070), .Q(
        interface3_bank_bus_dat_r[13]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[13]  ( .D(n3453), .CP(n6071), .Q(
        csrbank10_reload0_w[13]) );
  dfnrq1 \mgmtsoc_load_storage_reg[13]  ( .D(n3421), .CP(n6071), .Q(
        csrbank10_load0_w[13]) );
  dfnrq1 \mgmtsoc_value_reg[13]  ( .D(N5413), .CP(n6071), .Q(mgmtsoc_value[13]) );
  dfnrq1 \mgmtsoc_value_status_reg[13]  ( .D(n3487), .CP(n6071), .Q(
        csrbank10_value_w[13]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[13]  ( .D(N4707), .CP(n6071), .Q(
        interface10_bank_bus_dat_r[13]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[13]  ( .D(n3314), .CP(n6071), .Q(
        csrbank0_scratch0_w[13]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[13]  ( .D(N4112), .CP(n6071), .Q(
        interface0_bank_bus_dat_r[13]) );
  dfnrq1 \dbg_uart_data_reg[14]  ( .D(n3269), .CP(n6071), .Q(
        dbg_uart_wishbone_dat_w[14]) );
  dfnrq1 \la_out_storage_reg[14]  ( .D(n4466), .CP(n6072), .Q(n120) );
  dfnrq1 \la_out_storage_reg[46]  ( .D(n4434), .CP(n6072), .Q(n88) );
  dfnrq1 \la_out_storage_reg[78]  ( .D(n4402), .CP(n6072), .Q(n56) );
  dfnrq1 \la_out_storage_reg[110]  ( .D(n4370), .CP(n6072), .Q(n24) );
  dfnrq1 \la_oe_storage_reg[14]  ( .D(n4338), .CP(n6072), .Q(
        csrbank6_oe0_w[14]) );
  dfnrq1 \la_oe_storage_reg[46]  ( .D(n4306), .CP(n6072), .Q(
        csrbank6_oe1_w[14]) );
  dfnrq1 \la_oe_storage_reg[78]  ( .D(n4274), .CP(n6072), .Q(
        csrbank6_oe2_w[14]) );
  dfnrq1 \la_oe_storage_reg[110]  ( .D(n4242), .CP(n6072), .Q(
        csrbank6_oe3_w[14]) );
  dfnrq1 \la_ien_storage_reg[14]  ( .D(n4210), .CP(n6073), .Q(
        csrbank6_ien0_w[14]) );
  dfnrq1 \la_ien_storage_reg[46]  ( .D(n4178), .CP(n6073), .Q(
        csrbank6_ien1_w[14]) );
  dfnrq1 \la_ien_storage_reg[78]  ( .D(n4146), .CP(n6073), .Q(
        csrbank6_ien2_w[14]) );
  dfnrq1 \la_ien_storage_reg[110]  ( .D(n4114), .CP(n6073), .Q(
        csrbank6_ien3_w[14]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[14]  ( .D(N4477), .CP(n6073), .Q(
        interface6_bank_bus_dat_r[14]) );
  dfnrq1 \spimaster_storage_reg[14]  ( .D(n3706), .CP(n6073), .Q(
        spi_master_clk_divider0[14]) );
  dfnrq1 \spi_master_cs_storage_reg[14]  ( .D(n3667), .CP(n6073), .Q(
        csrbank9_cs0_w[14]) );
  dfnrq1 \spi_master_control_storage_reg[14]  ( .D(n3648), .CP(n6073), .Q(
        spi_master_length0[6]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[14]  ( .D(N4599), .CP(n6128), .Q(
        interface9_bank_bus_dat_r[14]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[14]  ( .D(n3588), 
        .CP(n6025), .Q(mgmtsoc_port_master_user_port_sink_payload_data[14]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[14]  ( .D(n3141), .CP(n6025), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[14]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[14]  ( .D(n3545), .CP(n6128), 
        .Q(csrbank3_master_phyconfig0_w[14]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[14]  ( .D(N4257), .CP(n6128), .Q(
        interface3_bank_bus_dat_r[14]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[14]  ( .D(n3452), .CP(n6025), .Q(
        csrbank10_reload0_w[14]) );
  dfnrq1 \mgmtsoc_load_storage_reg[14]  ( .D(n3420), .CP(n6128), .Q(
        csrbank10_load0_w[14]) );
  dfnrq1 \mgmtsoc_value_reg[14]  ( .D(N5414), .CP(n6025), .Q(mgmtsoc_value[14]) );
  dfnrq1 \mgmtsoc_value_status_reg[14]  ( .D(n3486), .CP(n6117), .Q(
        csrbank10_value_w[14]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[14]  ( .D(N4708), .CP(n6120), .Q(
        interface10_bank_bus_dat_r[14]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[14]  ( .D(n3313), .CP(n6068), .Q(
        csrbank0_scratch0_w[14]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[14]  ( .D(N4113), .CP(n6066), .Q(
        interface0_bank_bus_dat_r[14]) );
  dfnrq1 \dbg_uart_data_reg[15]  ( .D(n3268), .CP(n6117), .Q(
        dbg_uart_wishbone_dat_w[15]) );
  dfnrq1 \la_out_storage_reg[15]  ( .D(n4465), .CP(n6120), .Q(n119) );
  dfnrq1 \la_out_storage_reg[47]  ( .D(n4433), .CP(n6068), .Q(n87) );
  dfnrq1 \la_out_storage_reg[79]  ( .D(n4401), .CP(n6066), .Q(n55) );
  dfnrq1 \la_out_storage_reg[111]  ( .D(n4369), .CP(n6070), .Q(n23) );
  dfnrq1 \la_oe_storage_reg[15]  ( .D(n4337), .CP(n6071), .Q(
        csrbank6_oe0_w[15]) );
  dfnrq1 \la_oe_storage_reg[47]  ( .D(n4305), .CP(n6072), .Q(
        csrbank6_oe1_w[15]) );
  dfnrq1 \la_oe_storage_reg[79]  ( .D(n4273), .CP(n6073), .Q(
        csrbank6_oe2_w[15]) );
  dfnrq1 \la_oe_storage_reg[111]  ( .D(n4241), .CP(n6119), .Q(
        csrbank6_oe3_w[15]) );
  dfnrq1 \la_ien_storage_reg[15]  ( .D(n4209), .CP(n6070), .Q(
        csrbank6_ien0_w[15]) );
  dfnrq1 \la_ien_storage_reg[47]  ( .D(n4177), .CP(n6071), .Q(
        csrbank6_ien1_w[15]) );
  dfnrq1 \la_ien_storage_reg[79]  ( .D(n4145), .CP(n6024), .Q(
        csrbank6_ien2_w[15]) );
  dfnrq1 \la_ien_storage_reg[111]  ( .D(n4113), .CP(n6057), .Q(
        csrbank6_ien3_w[15]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[15]  ( .D(N4478), .CP(n6024), .Q(
        interface6_bank_bus_dat_r[15]) );
  dfnrq1 \spimaster_storage_reg[15]  ( .D(n3705), .CP(n6057), .Q(
        spi_master_clk_divider0[15]) );
  dfnrq1 \spi_master_cs_storage_reg[15]  ( .D(n3666), .CP(n6024), .Q(
        csrbank9_cs0_w[15]) );
  dfnrq1 \spi_master_control_storage_reg[15]  ( .D(n3647), .CP(n6057), .Q(
        spi_master_length0[7]) );
  dfnrq1 \interface9_bank_bus_dat_r_reg[15]  ( .D(N4600), .CP(n6024), .Q(
        interface9_bank_bus_dat_r[15]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[15]  ( .D(n3587), 
        .CP(n6057), .Q(mgmtsoc_port_master_user_port_sink_payload_data[15]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[15]  ( .D(n3142), .CP(n6074), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[15]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[16]  ( .D(n3143), .CP(n6074), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[16]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[15]  ( .D(n3544), .CP(n6074), 
        .Q(csrbank3_master_phyconfig0_w[15]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[15]  ( .D(N4258), .CP(n6074), .Q(
        interface3_bank_bus_dat_r[15]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[15]  ( .D(n3451), .CP(n6074), .Q(
        csrbank10_reload0_w[15]) );
  dfnrq1 \mgmtsoc_load_storage_reg[15]  ( .D(n3419), .CP(n6074), .Q(
        csrbank10_load0_w[15]) );
  dfnrq1 \mgmtsoc_value_reg[15]  ( .D(N5415), .CP(n6074), .Q(mgmtsoc_value[15]) );
  dfnrq1 \mgmtsoc_value_status_reg[15]  ( .D(n3485), .CP(n6074), .Q(
        csrbank10_value_w[15]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[15]  ( .D(N4709), .CP(n6075), .Q(
        interface10_bank_bus_dat_r[15]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[15]  ( .D(n3312), .CP(n6075), .Q(
        csrbank0_scratch0_w[15]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[15]  ( .D(N4114), .CP(n6075), .Q(
        interface0_bank_bus_dat_r[15]) );
  dfnrq1 \dbg_uart_data_reg[17]  ( .D(n3266), .CP(n6075), .Q(
        dbg_uart_wishbone_dat_w[17]) );
  dfnrq1 \la_out_storage_reg[17]  ( .D(n4463), .CP(n6075), .Q(n117) );
  dfnrq1 \la_out_storage_reg[49]  ( .D(n4431), .CP(n6075), .Q(n85) );
  dfnrq1 \la_out_storage_reg[81]  ( .D(n4399), .CP(n6075), .Q(n53) );
  dfnrq1 \la_out_storage_reg[113]  ( .D(n4367), .CP(n6075), .Q(n21) );
  dfnrq1 \la_oe_storage_reg[17]  ( .D(n4335), .CP(n6076), .Q(
        csrbank6_oe0_w[17]) );
  dfnrq1 \la_oe_storage_reg[49]  ( .D(n4303), .CP(n6076), .Q(
        csrbank6_oe1_w[17]) );
  dfnrq1 \la_oe_storage_reg[81]  ( .D(n4271), .CP(n6076), .Q(
        csrbank6_oe2_w[17]) );
  dfnrq1 \la_oe_storage_reg[113]  ( .D(n4239), .CP(n6076), .Q(
        csrbank6_oe3_w[17]) );
  dfnrq1 \la_ien_storage_reg[17]  ( .D(n4207), .CP(n6076), .Q(
        csrbank6_ien0_w[17]) );
  dfnrq1 \la_ien_storage_reg[49]  ( .D(n4175), .CP(n6076), .Q(
        csrbank6_ien1_w[17]) );
  dfnrq1 \la_ien_storage_reg[81]  ( .D(n4143), .CP(n6076), .Q(
        csrbank6_ien2_w[17]) );
  dfnrq1 \la_ien_storage_reg[113]  ( .D(n4111), .CP(n6076), .Q(
        csrbank6_ien3_w[17]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[17]  ( .D(N4480), .CP(n6077), .Q(
        interface6_bank_bus_dat_r[17]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[17]  ( .D(n3585), 
        .CP(n6077), .Q(mgmtsoc_port_master_user_port_sink_payload_data[17]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[17]  ( .D(n3144), .CP(n6077), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[17]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[17]  ( .D(n3542), .CP(n6077), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_mask[1]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[17]  ( .D(N4260), .CP(n6077), .Q(
        interface3_bank_bus_dat_r[17]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[17]  ( .D(n3449), .CP(n6077), .Q(
        csrbank10_reload0_w[17]) );
  dfnrq1 \mgmtsoc_load_storage_reg[17]  ( .D(n3417), .CP(n6077), .Q(
        csrbank10_load0_w[17]) );
  dfnrq1 \mgmtsoc_value_reg[17]  ( .D(N5417), .CP(n6077), .Q(mgmtsoc_value[17]) );
  dfnrq1 \mgmtsoc_value_status_reg[17]  ( .D(n3483), .CP(n6105), .Q(
        csrbank10_value_w[17]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[17]  ( .D(N4711), .CP(n6106), .Q(
        interface10_bank_bus_dat_r[17]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[17]  ( .D(n3310), .CP(n6104), .Q(
        csrbank0_scratch0_w[17]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[17]  ( .D(N4116), .CP(n6086), .Q(
        interface0_bank_bus_dat_r[17]) );
  dfnrq1 \dbg_uart_data_reg[18]  ( .D(n3265), .CP(n6123), .Q(
        dbg_uart_wishbone_dat_w[18]) );
  dfnrq1 \la_out_storage_reg[18]  ( .D(n4462), .CP(n6103), .Q(n116) );
  dfnrq1 \la_out_storage_reg[50]  ( .D(n4430), .CP(n6079), .Q(n84) );
  dfnrq1 \la_out_storage_reg[82]  ( .D(n4398), .CP(n6080), .Q(n52) );
  dfnrq1 \la_out_storage_reg[114]  ( .D(n4366), .CP(n6061), .Q(n20) );
  dfnrq1 \la_oe_storage_reg[18]  ( .D(n4334), .CP(n6081), .Q(
        csrbank6_oe0_w[18]) );
  dfnrq1 \la_oe_storage_reg[50]  ( .D(n4302), .CP(n6107), .Q(
        csrbank6_oe1_w[18]) );
  dfnrq1 \la_oe_storage_reg[82]  ( .D(n4270), .CP(n6090), .Q(
        csrbank6_oe2_w[18]) );
  dfnrq1 \la_oe_storage_reg[114]  ( .D(n4238), .CP(n6085), .Q(
        csrbank6_oe3_w[18]) );
  dfnrq1 \la_ien_storage_reg[18]  ( .D(n4206), .CP(n6074), .Q(
        csrbank6_ien0_w[18]) );
  dfnrq1 \la_ien_storage_reg[50]  ( .D(n4174), .CP(n6104), .Q(
        csrbank6_ien1_w[18]) );
  dfnrq1 \la_ien_storage_reg[82]  ( .D(n4142), .CP(n6075), .Q(
        csrbank6_ien2_w[18]) );
  dfnrq1 \la_ien_storage_reg[114]  ( .D(n4110), .CP(n6070), .Q(
        csrbank6_ien3_w[18]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[18]  ( .D(N4481), .CP(n6067), .Q(
        interface6_bank_bus_dat_r[18]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[18]  ( .D(n3584), 
        .CP(n6067), .Q(mgmtsoc_port_master_user_port_sink_payload_data[18]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[18]  ( .D(n3145), .CP(n6067), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[18]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[18]  ( .D(n3541), .CP(n6067), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_mask[2]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[18]  ( .D(N4261), .CP(n6067), .Q(
        interface3_bank_bus_dat_r[18]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[18]  ( .D(n3448), .CP(n6065), .Q(
        csrbank10_reload0_w[18]) );
  dfnrq1 \mgmtsoc_load_storage_reg[18]  ( .D(n3416), .CP(n6064), .Q(
        csrbank10_load0_w[18]) );
  dfnrq1 \mgmtsoc_value_reg[18]  ( .D(N5418), .CP(n6067), .Q(mgmtsoc_value[18]) );
  dfnrq1 \mgmtsoc_value_status_reg[18]  ( .D(n3482), .CP(n6067), .Q(
        csrbank10_value_w[18]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[18]  ( .D(N4712), .CP(n6119), .Q(
        interface10_bank_bus_dat_r[18]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[18]  ( .D(n3309), .CP(n6118), .Q(
        csrbank0_scratch0_w[18]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[18]  ( .D(N4117), .CP(n6065), .Q(
        interface0_bank_bus_dat_r[18]) );
  dfnrq1 \dbg_uart_data_reg[19]  ( .D(n3264), .CP(n6064), .Q(
        dbg_uart_wishbone_dat_w[19]) );
  dfnrq1 \la_out_storage_reg[19]  ( .D(n4461), .CP(n6065), .Q(n115) );
  dfnrq1 \la_out_storage_reg[51]  ( .D(n4429), .CP(n6064), .Q(n83) );
  dfnrq1 \la_out_storage_reg[83]  ( .D(n4397), .CP(n6067), .Q(n51) );
  dfnrq1 \la_out_storage_reg[115]  ( .D(n4365), .CP(n6064), .Q(n19) );
  dfnrq1 \la_oe_storage_reg[19]  ( .D(n4333), .CP(n6069), .Q(
        csrbank6_oe0_w[19]) );
  dfnrq1 \la_oe_storage_reg[51]  ( .D(n4301), .CP(n6065), .Q(
        csrbank6_oe1_w[19]) );
  dfnrq1 \la_oe_storage_reg[83]  ( .D(n4269), .CP(n6064), .Q(
        csrbank6_oe2_w[19]) );
  dfnrq1 \la_oe_storage_reg[115]  ( .D(n4237), .CP(n6067), .Q(
        csrbank6_oe3_w[19]) );
  dfnrq1 \la_ien_storage_reg[19]  ( .D(n4205), .CP(n6067), .Q(
        csrbank6_ien0_w[19]) );
  dfnrq1 \la_ien_storage_reg[51]  ( .D(n4173), .CP(n6118), .Q(
        csrbank6_ien1_w[19]) );
  dfnrq1 \la_ien_storage_reg[83]  ( .D(n4141), .CP(n6066), .Q(
        csrbank6_ien2_w[19]) );
  dfnrq1 \la_ien_storage_reg[115]  ( .D(n4109), .CP(n6065), .Q(
        csrbank6_ien3_w[19]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[19]  ( .D(N4482), .CP(n6064), .Q(
        interface6_bank_bus_dat_r[19]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[19]  ( .D(n3583), 
        .CP(n6067), .Q(mgmtsoc_port_master_user_port_sink_payload_data[19]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[19]  ( .D(n3146), .CP(n6118), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[19]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[19]  ( .D(n3540), .CP(n6068), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_mask[3]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[19]  ( .D(N4262), .CP(n6119), .Q(
        interface3_bank_bus_dat_r[19]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[19]  ( .D(n3447), .CP(n6119), .Q(
        csrbank10_reload0_w[19]) );
  dfnrq1 \mgmtsoc_load_storage_reg[19]  ( .D(n3415), .CP(n6070), .Q(
        csrbank10_load0_w[19]) );
  dfnrq1 \mgmtsoc_value_reg[19]  ( .D(N5419), .CP(n6071), .Q(mgmtsoc_value[19]) );
  dfnrq1 \mgmtsoc_value_status_reg[19]  ( .D(n3481), .CP(n6072), .Q(
        csrbank10_value_w[19]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[19]  ( .D(N4713), .CP(n6073), .Q(
        interface10_bank_bus_dat_r[19]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[19]  ( .D(n3308), .CP(n6069), .Q(
        csrbank0_scratch0_w[19]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[19]  ( .D(N4118), .CP(n6119), .Q(
        interface0_bank_bus_dat_r[19]) );
  dfnrq1 \dbg_uart_data_reg[20]  ( .D(n3263), .CP(n6073), .Q(
        dbg_uart_wishbone_dat_w[20]) );
  dfnrq1 \la_out_storage_reg[20]  ( .D(n4460), .CP(n6070), .Q(n114) );
  dfnrq1 \la_out_storage_reg[52]  ( .D(n4428), .CP(n6071), .Q(n82) );
  dfnrq1 \la_out_storage_reg[84]  ( .D(n4396), .CP(n6072), .Q(n50) );
  dfnrq1 \la_out_storage_reg[116]  ( .D(n4364), .CP(n6073), .Q(n18) );
  dfnrq1 \la_oe_storage_reg[20]  ( .D(n4332), .CP(n6069), .Q(
        csrbank6_oe0_w[20]) );
  dfnrq1 \la_oe_storage_reg[52]  ( .D(n4300), .CP(n6069), .Q(
        csrbank6_oe1_w[20]) );
  dfnrq1 \la_oe_storage_reg[84]  ( .D(n4268), .CP(n6119), .Q(
        csrbank6_oe2_w[20]) );
  dfnrq1 \la_oe_storage_reg[116]  ( .D(n4236), .CP(n6119), .Q(
        csrbank6_oe3_w[20]) );
  dfnrq1 \la_ien_storage_reg[20]  ( .D(n4204), .CP(n6069), .Q(
        csrbank6_ien0_w[20]) );
  dfnrq1 \la_ien_storage_reg[52]  ( .D(n4172), .CP(n6070), .Q(
        csrbank6_ien1_w[20]) );
  dfnrq1 \la_ien_storage_reg[84]  ( .D(n4140), .CP(n6071), .Q(
        csrbank6_ien2_w[20]) );
  dfnrq1 \la_ien_storage_reg[116]  ( .D(n4108), .CP(n6072), .Q(
        csrbank6_ien3_w[20]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[20]  ( .D(N4483), .CP(n6073), .Q(
        interface6_bank_bus_dat_r[20]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[20]  ( .D(n3582), 
        .CP(n6069), .Q(mgmtsoc_port_master_user_port_sink_payload_data[20]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[20]  ( .D(n3147), .CP(n6072), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[20]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[20]  ( .D(n3539), .CP(n6072), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_mask[4]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[20]  ( .D(N4263), .CP(n6073), .Q(
        interface3_bank_bus_dat_r[20]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[20]  ( .D(n3446), .CP(n6069), .Q(
        csrbank10_reload0_w[20]) );
  dfnrq1 \mgmtsoc_load_storage_reg[20]  ( .D(n3414), .CP(n6071), .Q(
        csrbank10_load0_w[20]) );
  dfnrq1 \mgmtsoc_value_reg[20]  ( .D(N5420), .CP(n6119), .Q(mgmtsoc_value[20]) );
  dfnrq1 \mgmtsoc_value_status_reg[20]  ( .D(n3480), .CP(n6071), .Q(
        csrbank10_value_w[20]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[20]  ( .D(N4714), .CP(n6072), .Q(
        interface10_bank_bus_dat_r[20]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[20]  ( .D(n3307), .CP(n6119), .Q(
        csrbank0_scratch0_w[20]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[20]  ( .D(N4119), .CP(n6119), .Q(
        interface0_bank_bus_dat_r[20]) );
  dfnrq1 \dbg_uart_data_reg[21]  ( .D(n3262), .CP(n6119), .Q(
        dbg_uart_wishbone_dat_w[21]) );
  dfnrq1 \la_out_storage_reg[21]  ( .D(n4459), .CP(n6073), .Q(n113) );
  dfnrq1 \la_out_storage_reg[53]  ( .D(n4427), .CP(n6070), .Q(n81) );
  dfnrq1 \la_out_storage_reg[85]  ( .D(n4395), .CP(n6071), .Q(n49) );
  dfnrq1 \la_out_storage_reg[117]  ( .D(n4363), .CP(n6072), .Q(n17) );
  dfnrq1 \la_oe_storage_reg[21]  ( .D(n4331), .CP(n6119), .Q(
        csrbank6_oe0_w[21]) );
  dfnrq1 \la_oe_storage_reg[53]  ( .D(n4299), .CP(n6068), .Q(
        csrbank6_oe1_w[21]) );
  dfnrq1 \la_oe_storage_reg[85]  ( .D(n4267), .CP(n6068), .Q(
        csrbank6_oe2_w[21]) );
  dfnrq1 \la_oe_storage_reg[117]  ( .D(n4235), .CP(n6068), .Q(
        csrbank6_oe3_w[21]) );
  dfnrq1 \la_ien_storage_reg[21]  ( .D(n4203), .CP(n6068), .Q(
        csrbank6_ien0_w[21]) );
  dfnrq1 \la_ien_storage_reg[53]  ( .D(n4171), .CP(n6068), .Q(
        csrbank6_ien1_w[21]) );
  dfnrq1 \la_ien_storage_reg[85]  ( .D(n4139), .CP(n6068), .Q(
        csrbank6_ien2_w[21]) );
  dfnrq1 \la_ien_storage_reg[117]  ( .D(n4107), .CP(n6068), .Q(
        csrbank6_ien3_w[21]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[21]  ( .D(N4484), .CP(n6068), .Q(
        interface6_bank_bus_dat_r[21]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[21]  ( .D(n3581), 
        .CP(n6069), .Q(mgmtsoc_port_master_user_port_sink_payload_data[21]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[21]  ( .D(n3148), .CP(n6069), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[21]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[21]  ( .D(n3538), .CP(n6069), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_mask[5]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[21]  ( .D(N4264), .CP(n6069), .Q(
        interface3_bank_bus_dat_r[21]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[21]  ( .D(n3445), .CP(n6069), .Q(
        csrbank10_reload0_w[21]) );
  dfnrq1 \mgmtsoc_load_storage_reg[21]  ( .D(n3413), .CP(n6069), .Q(
        csrbank10_load0_w[21]) );
  dfnrq1 \mgmtsoc_value_reg[21]  ( .D(N5421), .CP(n6069), .Q(mgmtsoc_value[21]) );
  dfnrq1 \mgmtsoc_value_status_reg[21]  ( .D(n3479), .CP(n6069), .Q(
        csrbank10_value_w[21]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[21]  ( .D(N4715), .CP(n6051), .Q(
        interface10_bank_bus_dat_r[21]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[21]  ( .D(n3306), .CP(n6098), .Q(
        csrbank0_scratch0_w[21]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[21]  ( .D(N4120), .CP(n6053), .Q(
        interface0_bank_bus_dat_r[21]) );
  dfnrq1 \dbg_uart_data_reg[22]  ( .D(n3261), .CP(n6055), .Q(
        dbg_uart_wishbone_dat_w[22]) );
  dfnrq1 \la_out_storage_reg[22]  ( .D(n4458), .CP(n6032), .Q(n112) );
  dfnrq1 \la_out_storage_reg[54]  ( .D(n4426), .CP(n6022), .Q(n80) );
  dfnrq1 \la_out_storage_reg[86]  ( .D(n4394), .CP(n6098), .Q(n48) );
  dfnrq1 \la_out_storage_reg[118]  ( .D(n4362), .CP(n6032), .Q(n16) );
  dfnrq1 \la_oe_storage_reg[22]  ( .D(n4330), .CP(n6118), .Q(
        csrbank6_oe0_w[22]) );
  dfnrq1 \la_oe_storage_reg[54]  ( .D(n4298), .CP(n6072), .Q(
        csrbank6_oe1_w[22]) );
  dfnrq1 \la_oe_storage_reg[86]  ( .D(n4266), .CP(n6118), .Q(
        csrbank6_oe2_w[22]) );
  dfnrq1 \la_oe_storage_reg[118]  ( .D(n4234), .CP(n6117), .Q(
        csrbank6_oe3_w[22]) );
  dfnrq1 \la_ien_storage_reg[22]  ( .D(n4202), .CP(n6120), .Q(
        csrbank6_ien0_w[22]) );
  dfnrq1 \la_ien_storage_reg[54]  ( .D(n4170), .CP(n6119), .Q(
        csrbank6_ien1_w[22]) );
  dfnrq1 \la_ien_storage_reg[86]  ( .D(n4138), .CP(n6065), .Q(
        csrbank6_ien2_w[22]) );
  dfnrq1 \la_ien_storage_reg[118]  ( .D(n4106), .CP(n6064), .Q(
        csrbank6_ien3_w[22]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[22]  ( .D(N4485), .CP(n6119), .Q(
        interface6_bank_bus_dat_r[22]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[22]  ( .D(n3580), 
        .CP(n6070), .Q(mgmtsoc_port_master_user_port_sink_payload_data[22]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[22]  ( .D(n3149), .CP(n6071), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[22]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[22]  ( .D(n3537), .CP(n6118), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_mask[6]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[22]  ( .D(N4265), .CP(n6117), .Q(
        interface3_bank_bus_dat_r[22]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[22]  ( .D(n3444), .CP(n6120), .Q(
        csrbank10_reload0_w[22]) );
  dfnrq1 \mgmtsoc_load_storage_reg[22]  ( .D(n3412), .CP(n6119), .Q(
        csrbank10_load0_w[22]) );
  dfnrq1 \mgmtsoc_value_reg[22]  ( .D(N5422), .CP(n6072), .Q(mgmtsoc_value[22]) );
  dfnrq1 \mgmtsoc_value_status_reg[22]  ( .D(n3478), .CP(n6069), .Q(
        csrbank10_value_w[22]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[22]  ( .D(N4716), .CP(n6119), .Q(
        interface10_bank_bus_dat_r[22]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[22]  ( .D(n3305), .CP(n6063), .Q(
        csrbank0_scratch0_w[22]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[22]  ( .D(N4121), .CP(n6073), .Q(
        interface0_bank_bus_dat_r[22]) );
  dfnrq1 \dbg_uart_data_reg[23]  ( .D(n3260), .CP(n6117), .Q(
        dbg_uart_wishbone_dat_w[23]) );
  dfnrq1 \la_out_storage_reg[23]  ( .D(n4457), .CP(n6120), .Q(n111) );
  dfnrq1 \la_out_storage_reg[55]  ( .D(n4425), .CP(n6118), .Q(n79) );
  dfnrq1 \la_out_storage_reg[87]  ( .D(n4393), .CP(n6069), .Q(n47) );
  dfnrq1 \la_out_storage_reg[119]  ( .D(n4361), .CP(n6073), .Q(n15) );
  dfnrq1 \la_oe_storage_reg[23]  ( .D(n4329), .CP(n6066), .Q(
        csrbank6_oe0_w[23]) );
  dfnrq1 \la_oe_storage_reg[55]  ( .D(n4297), .CP(n6122), .Q(
        csrbank6_oe1_w[23]) );
  dfnrq1 \la_oe_storage_reg[87]  ( .D(n4265), .CP(n6084), .Q(
        csrbank6_oe2_w[23]) );
  dfnrq1 \la_oe_storage_reg[119]  ( .D(n4233), .CP(n6084), .Q(
        csrbank6_oe3_w[23]) );
  dfnrq1 \la_ien_storage_reg[23]  ( .D(n4201), .CP(n6061), .Q(
        csrbank6_ien0_w[23]) );
  dfnrq1 \la_ien_storage_reg[55]  ( .D(n4169), .CP(n6084), .Q(
        csrbank6_ien1_w[23]) );
  dfnrq1 \la_ien_storage_reg[87]  ( .D(n4137), .CP(n6084), .Q(
        csrbank6_ien2_w[23]) );
  dfnrq1 \la_ien_storage_reg[119]  ( .D(n4105), .CP(n6084), .Q(
        csrbank6_ien3_w[23]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[23]  ( .D(N4486), .CP(n6084), .Q(
        interface6_bank_bus_dat_r[23]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[23]  ( .D(n3579), 
        .CP(n6084), .Q(mgmtsoc_port_master_user_port_sink_payload_data[23]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[23]  ( .D(n3150), .CP(n6084), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[23]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[24]  ( .D(n3151), .CP(n6085), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[24]) );
  dfnrq1 \mgmtsoc_master_phyconfig_storage_reg[23]  ( .D(n3536), .CP(n6085), 
        .Q(mgmtsoc_master_tx_fifo_sink_payload_mask[7]) );
  dfnrq1 \interface3_bank_bus_dat_r_reg[23]  ( .D(N4266), .CP(n6085), .Q(
        interface3_bank_bus_dat_r[23]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[23]  ( .D(n3443), .CP(n6085), .Q(
        csrbank10_reload0_w[23]) );
  dfnrq1 \mgmtsoc_load_storage_reg[23]  ( .D(n3411), .CP(n6085), .Q(
        csrbank10_load0_w[23]) );
  dfnrq1 \mgmtsoc_value_reg[23]  ( .D(N5423), .CP(n6085), .Q(mgmtsoc_value[23]) );
  dfnrq1 \mgmtsoc_value_status_reg[23]  ( .D(n3477), .CP(n6085), .Q(
        csrbank10_value_w[23]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[23]  ( .D(N4717), .CP(n6085), .Q(
        interface10_bank_bus_dat_r[23]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[23]  ( .D(n3304), .CP(n6086), .Q(
        csrbank0_scratch0_w[23]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[23]  ( .D(N4122), .CP(n6086), .Q(
        interface0_bank_bus_dat_r[23]) );
  dfnrq1 \dbg_uart_data_reg[25]  ( .D(n3258), .CP(n6086), .Q(
        dbg_uart_wishbone_dat_w[25]) );
  dfnrq1 \la_out_storage_reg[25]  ( .D(n4455), .CP(n6086), .Q(n109) );
  dfnrq1 \la_out_storage_reg[57]  ( .D(n4423), .CP(n6086), .Q(n77) );
  dfnrq1 \la_out_storage_reg[89]  ( .D(n4391), .CP(n6086), .Q(n45) );
  dfnrq1 \la_out_storage_reg[121]  ( .D(n4359), .CP(n6086), .Q(n13) );
  dfnrq1 \la_oe_storage_reg[25]  ( .D(n4327), .CP(n6086), .Q(
        csrbank6_oe0_w[25]) );
  dfnrq1 \la_oe_storage_reg[57]  ( .D(n4295), .CP(n6123), .Q(
        csrbank6_oe1_w[25]) );
  dfnrq1 \la_oe_storage_reg[89]  ( .D(n4263), .CP(n6123), .Q(
        csrbank6_oe2_w[25]) );
  dfnrq1 \la_oe_storage_reg[121]  ( .D(n4231), .CP(n6101), .Q(
        csrbank6_oe3_w[25]) );
  dfnrq1 \la_ien_storage_reg[25]  ( .D(n4199), .CP(n6079), .Q(
        csrbank6_ien0_w[25]) );
  dfnrq1 \la_ien_storage_reg[57]  ( .D(n4167), .CP(n6074), .Q(
        csrbank6_ien1_w[25]) );
  dfnrq1 \la_ien_storage_reg[89]  ( .D(n4135), .CP(n6075), .Q(
        csrbank6_ien2_w[25]) );
  dfnrq1 \la_ien_storage_reg[121]  ( .D(n4103), .CP(n6124), .Q(
        csrbank6_ien3_w[25]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[25]  ( .D(N4488), .CP(n6079), .Q(
        interface6_bank_bus_dat_r[25]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[25]  ( .D(n3577), 
        .CP(n6096), .Q(mgmtsoc_port_master_user_port_sink_payload_data[25]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[25]  ( .D(n3152), .CP(n6085), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[25]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[25]  ( .D(n3441), .CP(n6079), .Q(
        csrbank10_reload0_w[25]) );
  dfnrq1 \mgmtsoc_load_storage_reg[25]  ( .D(n3409), .CP(n6076), .Q(
        csrbank10_load0_w[25]) );
  dfnrq1 \mgmtsoc_value_reg[25]  ( .D(N5425), .CP(n6033), .Q(mgmtsoc_value[25]) );
  dfnrq1 \mgmtsoc_value_status_reg[25]  ( .D(n3475), .CP(n6077), .Q(
        csrbank10_value_w[25]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[25]  ( .D(N4719), .CP(n6123), .Q(
        interface10_bank_bus_dat_r[25]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[25]  ( .D(n3302), .CP(n6079), .Q(
        csrbank0_scratch0_w[25]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[25]  ( .D(N4124), .CP(n6128), .Q(
        interface0_bank_bus_dat_r[25]) );
  dfnrq1 \dbg_uart_data_reg[26]  ( .D(n3257), .CP(n6123), .Q(
        dbg_uart_wishbone_dat_w[26]) );
  dfnrq1 \la_out_storage_reg[26]  ( .D(n4454), .CP(n6123), .Q(n108) );
  dfnrq1 \la_out_storage_reg[58]  ( .D(n4422), .CP(n6079), .Q(n76) );
  dfnrq1 \la_out_storage_reg[90]  ( .D(n4390), .CP(n6042), .Q(n44) );
  dfnrq1 \la_out_storage_reg[122]  ( .D(n4358), .CP(n6082), .Q(n12) );
  dfnrq1 \la_oe_storage_reg[26]  ( .D(n4326), .CP(n6082), .Q(
        csrbank6_oe0_w[26]) );
  dfnrq1 \la_oe_storage_reg[58]  ( .D(n4294), .CP(n6033), .Q(
        csrbank6_oe1_w[26]) );
  dfnrq1 \la_oe_storage_reg[90]  ( .D(n4262), .CP(n6081), .Q(
        csrbank6_oe2_w[26]) );
  dfnrq1 \la_oe_storage_reg[122]  ( .D(n4230), .CP(n6079), .Q(
        csrbank6_oe3_w[26]) );
  dfnrq1 \la_ien_storage_reg[26]  ( .D(n4198), .CP(n6033), .Q(
        csrbank6_ien0_w[26]) );
  dfnrq1 \la_ien_storage_reg[58]  ( .D(n4166), .CP(n6123), .Q(
        csrbank6_ien1_w[26]) );
  dfnrq1 \la_ien_storage_reg[90]  ( .D(n4134), .CP(n6043), .Q(
        csrbank6_ien2_w[26]) );
  dfnrq1 \la_ien_storage_reg[122]  ( .D(n4102), .CP(n6080), .Q(
        csrbank6_ien3_w[26]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[26]  ( .D(N4489), .CP(n6082), .Q(
        interface6_bank_bus_dat_r[26]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[26]  ( .D(n3576), 
        .CP(n6123), .Q(mgmtsoc_port_master_user_port_sink_payload_data[26]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[26]  ( .D(n3153), .CP(n6122), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[26]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[26]  ( .D(n3440), .CP(n6122), .Q(
        csrbank10_reload0_w[26]) );
  dfnrq1 \mgmtsoc_load_storage_reg[26]  ( .D(n3408), .CP(n6121), .Q(
        csrbank10_load0_w[26]) );
  dfnrq1 \mgmtsoc_value_reg[26]  ( .D(N5426), .CP(n6121), .Q(mgmtsoc_value[26]) );
  dfnrq1 \mgmtsoc_value_status_reg[26]  ( .D(n3474), .CP(n6121), .Q(
        csrbank10_value_w[26]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[26]  ( .D(N4720), .CP(n6122), .Q(
        interface10_bank_bus_dat_r[26]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[26]  ( .D(n3301), .CP(n6122), .Q(
        csrbank0_scratch0_w[26]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[26]  ( .D(N4125), .CP(n6086), .Q(
        interface0_bank_bus_dat_r[26]) );
  dfnrq1 \dbg_uart_data_reg[27]  ( .D(n3256), .CP(n6122), .Q(
        dbg_uart_wishbone_dat_w[27]) );
  dfnrq1 \la_out_storage_reg[27]  ( .D(n4453), .CP(n6122), .Q(n107) );
  dfnrq1 \la_out_storage_reg[59]  ( .D(n4421), .CP(n6121), .Q(n75) );
  dfnrq1 \la_out_storage_reg[91]  ( .D(n4389), .CP(n6122), .Q(n43) );
  dfnrq1 \la_out_storage_reg[123]  ( .D(n4357), .CP(n6121), .Q(n11) );
  dfnrq1 \la_oe_storage_reg[27]  ( .D(n4325), .CP(n6121), .Q(
        csrbank6_oe0_w[27]) );
  dfnrq1 \la_oe_storage_reg[59]  ( .D(n4293), .CP(n6122), .Q(
        csrbank6_oe1_w[27]) );
  dfnrq1 \la_oe_storage_reg[91]  ( .D(n4261), .CP(n6122), .Q(
        csrbank6_oe2_w[27]) );
  dfnrq1 \la_oe_storage_reg[123]  ( .D(n4229), .CP(n6121), .Q(
        csrbank6_oe3_w[27]) );
  dfnrq1 \la_ien_storage_reg[27]  ( .D(n4197), .CP(n6121), .Q(
        csrbank6_ien0_w[27]) );
  dfnrq1 \la_ien_storage_reg[59]  ( .D(n4165), .CP(n6122), .Q(
        csrbank6_ien1_w[27]) );
  dfnrq1 \la_ien_storage_reg[91]  ( .D(n4133), .CP(n6083), .Q(
        csrbank6_ien2_w[27]) );
  dfnrq1 \la_ien_storage_reg[123]  ( .D(n4101), .CP(n6084), .Q(
        csrbank6_ien3_w[27]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[27]  ( .D(N4490), .CP(n6085), .Q(
        interface6_bank_bus_dat_r[27]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[27]  ( .D(n3575), 
        .CP(n6122), .Q(mgmtsoc_port_master_user_port_sink_payload_data[27]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[27]  ( .D(n3154), .CP(n6086), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[27]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[27]  ( .D(n3439), .CP(n6122), .Q(
        csrbank10_reload0_w[27]) );
  dfnrq1 \mgmtsoc_load_storage_reg[27]  ( .D(n3407), .CP(n6122), .Q(
        csrbank10_load0_w[27]) );
  dfnrq1 \mgmtsoc_value_reg[27]  ( .D(N5427), .CP(n6121), .Q(mgmtsoc_value[27]) );
  dfnrq1 \mgmtsoc_value_status_reg[27]  ( .D(n3473), .CP(n6083), .Q(
        csrbank10_value_w[27]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[27]  ( .D(N4721), .CP(n6084), .Q(
        interface10_bank_bus_dat_r[27]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[27]  ( .D(n3300), .CP(n6085), .Q(
        csrbank0_scratch0_w[27]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[27]  ( .D(N4126), .CP(n6086), .Q(
        interface0_bank_bus_dat_r[27]) );
  dfnrq1 \la_out_storage_reg[28]  ( .D(n4452), .CP(n6100), .Q(n106) );
  dfnrq1 \la_out_storage_reg[60]  ( .D(n4420), .CP(n6085), .Q(n74) );
  dfnrq1 \la_out_storage_reg[92]  ( .D(n4388), .CP(n6105), .Q(n42) );
  dfnrq1 \la_out_storage_reg[124]  ( .D(n4356), .CP(n6033), .Q(n10) );
  dfnrq1 \la_oe_storage_reg[28]  ( .D(n4324), .CP(n6086), .Q(
        csrbank6_oe0_w[28]) );
  dfnrq1 \la_oe_storage_reg[60]  ( .D(n4292), .CP(n6078), .Q(
        csrbank6_oe1_w[28]) );
  dfnrq1 \la_oe_storage_reg[92]  ( .D(n4260), .CP(n6113), .Q(
        csrbank6_oe2_w[28]) );
  dfnrq1 \la_oe_storage_reg[124]  ( .D(n4228), .CP(n6085), .Q(
        csrbank6_oe3_w[28]) );
  dfnrq1 \la_ien_storage_reg[28]  ( .D(n4196), .CP(n6082), .Q(
        csrbank6_ien0_w[28]) );
  dfnrq1 \la_ien_storage_reg[60]  ( .D(n4164), .CP(n6033), .Q(
        csrbank6_ien1_w[28]) );
  dfnrq1 \la_ien_storage_reg[92]  ( .D(n4132), .CP(n6086), .Q(
        csrbank6_ien2_w[28]) );
  dfnrq1 \la_ien_storage_reg[124]  ( .D(n4100), .CP(n6116), .Q(
        csrbank6_ien3_w[28]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[28]  ( .D(N4491), .CP(n6097), .Q(
        interface6_bank_bus_dat_r[28]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[28]  ( .D(n3574), 
        .CP(n6076), .Q(mgmtsoc_port_master_user_port_sink_payload_data[28]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[28]  ( .D(n3155), .CP(n6085), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[28]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[28]  ( .D(n3438), .CP(n6086), .Q(
        csrbank10_reload0_w[28]) );
  dfnrq1 \mgmtsoc_load_storage_reg[28]  ( .D(n3406), .CP(n6082), .Q(
        csrbank10_load0_w[28]) );
  dfnrq1 \mgmtsoc_value_reg[28]  ( .D(N5428), .CP(n6080), .Q(mgmtsoc_value[28]) );
  dfnrq1 \mgmtsoc_value_status_reg[28]  ( .D(n3472), .CP(n6123), .Q(
        csrbank10_value_w[28]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[28]  ( .D(N4722), .CP(n6033), .Q(
        interface10_bank_bus_dat_r[28]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[28]  ( .D(n3299), .CP(n6090), .Q(
        csrbank0_scratch0_w[28]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[28]  ( .D(N4127), .CP(n6092), .Q(
        interface0_bank_bus_dat_r[28]) );
  dfnrq1 \la_out_storage_reg[29]  ( .D(n4451), .CP(n6093), .Q(n105) );
  dfnrq1 \la_out_storage_reg[61]  ( .D(n4419), .CP(n6096), .Q(n73) );
  dfnrq1 \la_out_storage_reg[93]  ( .D(n4387), .CP(n6123), .Q(n41) );
  dfnrq1 \la_out_storage_reg[125]  ( .D(n4355), .CP(n6097), .Q(n9) );
  dfnrq1 \la_oe_storage_reg[29]  ( .D(n4323), .CP(n6076), .Q(
        csrbank6_oe0_w[29]) );
  dfnrq1 \la_oe_storage_reg[61]  ( .D(n4291), .CP(n6089), .Q(
        csrbank6_oe1_w[29]) );
  dfnrq1 \la_oe_storage_reg[93]  ( .D(n4259), .CP(n6024), .Q(
        csrbank6_oe2_w[29]) );
  dfnrq1 \la_oe_storage_reg[125]  ( .D(n4227), .CP(n6054), .Q(
        csrbank6_oe3_w[29]) );
  dfnrq1 \la_ien_storage_reg[29]  ( .D(n4195), .CP(n6059), .Q(
        csrbank6_ien0_w[29]) );
  dfnrq1 \la_ien_storage_reg[61]  ( .D(n4163), .CP(n6080), .Q(
        csrbank6_ien1_w[29]) );
  dfnrq1 \la_ien_storage_reg[93]  ( .D(n4131), .CP(n6081), .Q(
        csrbank6_ien2_w[29]) );
  dfnrq1 \la_ien_storage_reg[125]  ( .D(n4099), .CP(n6105), .Q(
        csrbank6_ien3_w[29]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[29]  ( .D(N4492), .CP(n6094), .Q(
        interface6_bank_bus_dat_r[29]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[29]  ( .D(n3573), 
        .CP(n6106), .Q(mgmtsoc_port_master_user_port_sink_payload_data[29]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[29]  ( .D(n3156), .CP(n6048), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[29]) );
  dfnrq1 \mgmtsoc_reload_storage_reg[29]  ( .D(n3437), .CP(n6129), .Q(
        csrbank10_reload0_w[29]) );
  dfnrq1 \mgmtsoc_load_storage_reg[29]  ( .D(n3405), .CP(n6041), .Q(
        csrbank10_load0_w[29]) );
  dfnrq1 \mgmtsoc_value_reg[29]  ( .D(N5429), .CP(n6109), .Q(mgmtsoc_value[29]) );
  dfnrq1 \mgmtsoc_value_status_reg[29]  ( .D(n3471), .CP(n6110), .Q(
        csrbank10_value_w[29]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[29]  ( .D(N4723), .CP(n6080), .Q(
        interface10_bank_bus_dat_r[29]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[29]  ( .D(n3298), .CP(n6054), .Q(
        csrbank0_scratch0_w[29]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[29]  ( .D(N4128), .CP(n6079), .Q(
        interface0_bank_bus_dat_r[29]) );
  dfnrq1 \la_out_storage_reg[30]  ( .D(n4450), .CP(n6077), .Q(n104) );
  dfnrq1 \la_out_storage_reg[62]  ( .D(n4418), .CP(n6109), .Q(n72) );
  dfnrq1 \la_out_storage_reg[94]  ( .D(n4386), .CP(n6076), .Q(n40) );
  dfnrq1 \la_out_storage_reg[126]  ( .D(n4354), .CP(n6078), .Q(n8) );
  dfnrq1 \la_oe_storage_reg[30]  ( .D(n4322), .CP(n6078), .Q(
        csrbank6_oe0_w[30]) );
  dfnrq1 \la_oe_storage_reg[62]  ( .D(n4290), .CP(n6078), .Q(
        csrbank6_oe1_w[30]) );
  dfnrq1 \la_oe_storage_reg[94]  ( .D(n4258), .CP(n6078), .Q(
        csrbank6_oe2_w[30]) );
  dfnrq1 \la_oe_storage_reg[126]  ( .D(n4226), .CP(n6078), .Q(
        csrbank6_oe3_w[30]) );
  dfnrq1 \la_ien_storage_reg[30]  ( .D(n4194), .CP(n6078), .Q(
        csrbank6_ien0_w[30]) );
  dfnrq1 \la_ien_storage_reg[62]  ( .D(n4162), .CP(n6078), .Q(
        csrbank6_ien1_w[30]) );
  dfnrq1 \la_ien_storage_reg[94]  ( .D(n4130), .CP(n6078), .Q(
        csrbank6_ien2_w[30]) );
  dfnrq1 \la_ien_storage_reg[126]  ( .D(n4098), .CP(n6079), .Q(
        csrbank6_ien3_w[30]) );
  dfnrq1 \interface6_bank_bus_dat_r_reg[30]  ( .D(N4493), .CP(n6078), .Q(
        interface6_bank_bus_dat_r[30]) );
  dfnrq1 \mgmtsoc_master_tx_fifo_source_payload_data_reg[30]  ( .D(n3572), 
        .CP(n6080), .Q(mgmtsoc_port_master_user_port_sink_payload_data[30]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[30]  ( .D(n3157), .CP(n6081), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[30]) );
  dfnrq1 \mgmtsoc_litespisdrphycore_sr_out_reg[31]  ( .D(n3158), .CP(n6092), 
        .Q(mgmtsoc_litespisdrphycore_sr_out[31]) );
  dfnrq1 flash_io0_do_reg ( .D(mgmtsoc_litespisdrphycore_dq_o), .CP(n6123), 
        .Q(flash_io0_do) );
  dfnrq1 \mgmtsoc_reload_storage_reg[30]  ( .D(n3436), .CP(n6082), .Q(
        csrbank10_reload0_w[30]) );
  dfnrq1 \mgmtsoc_load_storage_reg[30]  ( .D(n3404), .CP(n6082), .Q(
        csrbank10_load0_w[30]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[30]  ( .D(n3297), .CP(n6102), .Q(
        csrbank0_scratch0_w[30]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[30]  ( .D(N4129), .CP(n6074), .Q(
        interface0_bank_bus_dat_r[30]) );
  dfnrq1 mgmtsoc_zero_pending_reg ( .D(n3501), .CP(n6078), .Q(mgmtsoc_zero1)
         );
  dfnrq1 \interface10_bank_bus_dat_r_reg[0]  ( .D(N4694), .CP(n6075), .Q(
        interface10_bank_bus_dat_r[0]) );
  dfnrq1 \mgmtsoc_value_status_reg[31]  ( .D(n3469), .CP(n6078), .Q(
        csrbank10_value_w[31]) );
  dfnrq1 \interface10_bank_bus_dat_r_reg[31]  ( .D(N4725), .CP(n6078), .Q(
        interface10_bank_bus_dat_r[31]) );
  dfnrq1 \mgmtsoc_scratch_storage_reg[31]  ( .D(n3296), .CP(n6076), .Q(
        csrbank0_scratch0_w[31]) );
  dfnrq1 \interface0_bank_bus_dat_r_reg[31]  ( .D(N4130), .CP(n6077), .Q(
        interface0_bank_bus_dat_r[31]) );
  dfnrq1 \dbg_uart_tx_data_reg[7]  ( .D(n3088), .CP(n6078), .Q(
        dbg_uart_tx_data[7]) );
  dfnrq1 \dbg_uart_tx_data_reg[6]  ( .D(n3090), .CP(n6083), .Q(
        dbg_uart_tx_data[6]) );
  dfnrq1 \dbg_uart_tx_data_reg[5]  ( .D(n3091), .CP(n6078), .Q(
        dbg_uart_tx_data[5]) );
  dfnrq1 \dbg_uart_tx_data_reg[4]  ( .D(n3092), .CP(n6085), .Q(
        dbg_uart_tx_data[4]) );
  dfnrq1 \dbg_uart_tx_data_reg[3]  ( .D(n3093), .CP(n6078), .Q(
        dbg_uart_tx_data[3]) );
  dfnrq1 \dbg_uart_tx_data_reg[2]  ( .D(n3094), .CP(n6084), .Q(
        dbg_uart_tx_data[2]) );
  dfnrq1 \dbg_uart_tx_data_reg[1]  ( .D(n3095), .CP(n6078), .Q(
        dbg_uart_tx_data[1]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[0]  ( .D(n3221), .CP(n6033), .Q(
        mgmtsoc_litespimmap_burst_adr[0]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[1]  ( .D(n3220), .CP(n6079), .Q(
        mgmtsoc_litespimmap_burst_adr[1]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[2]  ( .D(n3219), .CP(n6079), .Q(
        mgmtsoc_litespimmap_burst_adr[2]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[3]  ( .D(n3218), .CP(n6079), .Q(
        mgmtsoc_litespimmap_burst_adr[3]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[4]  ( .D(n3217), .CP(n6079), .Q(
        mgmtsoc_litespimmap_burst_adr[4]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[5]  ( .D(n3216), .CP(n6079), .Q(
        mgmtsoc_litespimmap_burst_adr[5]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[6]  ( .D(n3215), .CP(n6079), .Q(
        mgmtsoc_litespimmap_burst_adr[6]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[7]  ( .D(n3214), .CP(n6079), .Q(
        mgmtsoc_litespimmap_burst_adr[7]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[8]  ( .D(n3213), .CP(n6079), .Q(
        mgmtsoc_litespimmap_burst_adr[8]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[9]  ( .D(n3212), .CP(n6080), .Q(
        mgmtsoc_litespimmap_burst_adr[9]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[10]  ( .D(n3211), .CP(n6080), .Q(
        mgmtsoc_litespimmap_burst_adr[10]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[11]  ( .D(n3210), .CP(n6080), .Q(
        mgmtsoc_litespimmap_burst_adr[11]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[12]  ( .D(n3209), .CP(n6080), .Q(
        mgmtsoc_litespimmap_burst_adr[12]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[13]  ( .D(n3208), .CP(n6080), .Q(
        mgmtsoc_litespimmap_burst_adr[13]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[14]  ( .D(n3207), .CP(n6080), .Q(
        mgmtsoc_litespimmap_burst_adr[14]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[15]  ( .D(n3206), .CP(n6080), .Q(
        mgmtsoc_litespimmap_burst_adr[15]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[16]  ( .D(n3205), .CP(n6081), .Q(
        mgmtsoc_litespimmap_burst_adr[16]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[17]  ( .D(n3204), .CP(n6081), .Q(
        mgmtsoc_litespimmap_burst_adr[17]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[18]  ( .D(n3203), .CP(n6081), .Q(
        mgmtsoc_litespimmap_burst_adr[18]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[19]  ( .D(n3202), .CP(n6081), .Q(
        mgmtsoc_litespimmap_burst_adr[19]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[20]  ( .D(n3201), .CP(n6081), .Q(
        mgmtsoc_litespimmap_burst_adr[20]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[21]  ( .D(n3200), .CP(n6081), .Q(
        mgmtsoc_litespimmap_burst_adr[21]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[22]  ( .D(n3199), .CP(n6081), .Q(
        mgmtsoc_litespimmap_burst_adr[22]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[23]  ( .D(n3198), .CP(n6081), .Q(
        mgmtsoc_litespimmap_burst_adr[23]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[24]  ( .D(n3197), .CP(n6039), .Q(
        mgmtsoc_litespimmap_burst_adr[24]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[25]  ( .D(n3196), .CP(n6026), .Q(
        mgmtsoc_litespimmap_burst_adr[25]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[26]  ( .D(n3195), .CP(n6029), .Q(
        mgmtsoc_litespimmap_burst_adr[26]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[27]  ( .D(n3194), .CP(n6057), .Q(
        mgmtsoc_litespimmap_burst_adr[27]) );
  dfnrq1 \mgmtsoc_litespimmap_burst_adr_reg[28]  ( .D(n3193), .CP(n6056), .Q(
        mgmtsoc_litespimmap_burst_adr[28]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[0]  ( .D(n3399), .CP(n6091), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[0]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[1]  ( .D(n3398), .CP(n6121), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[1]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[2]  ( .D(n3397), .CP(n6105), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[2]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[3]  ( .D(n3396), .CP(n6082), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[3]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[4]  ( .D(n3395), .CP(n6080), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[4]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[5]  ( .D(n3394), .CP(n6081), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[5]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[6]  ( .D(n3393), .CP(n6045), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[6]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[7]  ( .D(n3392), .CP(n6044), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[7]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[8]  ( .D(n3391), .CP(n6049), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[8]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[9]  ( .D(n3390), .CP(n6123), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[9]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[10]  ( .D(n3389), .CP(n6080), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[10]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[11]  ( .D(n3388), .CP(n6033), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[11]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[12]  ( .D(n3387), .CP(n6080), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[12]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[13]  ( .D(n3386), .CP(n6086), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[13]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[14]  ( .D(n3385), .CP(n6080), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[14]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[15]  ( .D(n3384), .CP(n6082), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[15]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[16]  ( .D(n3383), .CP(n6080), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[16]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[17]  ( .D(n3382), .CP(n6082), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[17]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[18]  ( .D(n3381), .CP(n6082), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[18]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[19]  ( .D(n3380), .CP(n6082), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[19]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[20]  ( .D(n3379), .CP(n6082), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[20]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[21]  ( .D(n3378), .CP(n6082), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[21]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[22]  ( .D(n3377), .CP(n6082), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[22]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[23]  ( .D(n3376), .CP(n6082), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[23]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[24]  ( .D(n3375), .CP(n6082), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[24]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[25]  ( .D(n3374), .CP(n6125), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[25]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[26]  ( .D(n3373), .CP(n6081), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[26]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[27]  ( .D(n3372), .CP(n6097), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[27]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[28]  ( .D(n3371), .CP(n6081), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[28]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[29]  ( .D(n3370), .CP(n6076), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[29]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[30]  ( .D(n3369), .CP(n6081), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[30]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_data_reg[31]  ( .D(n3368), .CP(n6085), 
        .Q(mgmtsoc_vexriscv_i_cmd_payload_data[31]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_address_reg[2]  ( .D(n3367), .CP(
        n6081), .Q(mgmtsoc_vexriscv_i_cmd_payload_address[2]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_address_reg[3]  ( .D(n3366), .CP(
        n6083), .Q(mgmtsoc_vexriscv_i_cmd_payload_address[3]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_address_reg[4]  ( .D(n3365), .CP(
        n6083), .Q(mgmtsoc_vexriscv_i_cmd_payload_address[4]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_address_reg[5]  ( .D(n3364), .CP(
        n6083), .Q(mgmtsoc_vexriscv_i_cmd_payload_address[5]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_address_reg[6]  ( .D(n3363), .CP(
        n6083), .Q(mgmtsoc_vexriscv_i_cmd_payload_address[6]) );
  dfnrq1 \mgmtsoc_vexriscv_i_cmd_payload_address_reg[7]  ( .D(n3362), .CP(
        n6083), .Q(mgmtsoc_vexriscv_i_cmd_payload_address[7]) );
  dfnrq1 mgmtsoc_vexriscv_i_cmd_payload_wr_reg ( .D(n3361), .CP(n6083), .Q(
        mgmtsoc_vexriscv_i_cmd_payload_wr) );
  dfnrq1 \dbg_uart_tx_data_reg[0]  ( .D(n3096), .CP(n6083), .Q(
        dbg_uart_tx_data[0]) );
  dfnrq1 dbg_uart_dbg_uart_tx_reg ( .D(n4067), .CP(n6083), .Q(
        dbg_uart_dbg_uart_tx) );
  dfnrq1 \spimaster_storage_reg[0]  ( .D(n3720), .CP(n6058), .Q(
        spi_master_clk_divider0[0]) );
  dfnrq1 \spimaster_storage_reg[2]  ( .D(n3718), .CP(n6088), .Q(
        spi_master_clk_divider0[2]) );
  or02d4 U3 ( .A1(n2300), .A2(n5111), .Z(n2328) );
  inv0d1 U4 ( .I(uart_phy_rx_data[6]), .ZN(n3053) );
  inv0d1 U5 ( .I(uart_phy_rx_data[4]), .ZN(n3051) );
  inv0d1 U6 ( .I(n5990), .ZN(n5987) );
  nd02d1 U7 ( .A1(n4580), .A2(n4579), .ZN(n4581) );
  inv0d1 U8 ( .I(n5862), .ZN(n5830) );
  inv0d1 U9 ( .I(n5111), .ZN(n5340) );
  inv0d0 U10 ( .I(n4582), .ZN(n266) );
  nd04d0 U11 ( .A1(n760), .A2(n759), .A3(n758), .A4(n757), .ZN(N4480) );
  nd04d0 U12 ( .A1(n831), .A2(n830), .A3(n829), .A4(n828), .ZN(N4484) );
  nd04d0 U13 ( .A1(n889), .A2(n888), .A3(n887), .A4(n886), .ZN(N4486) );
  nd04d0 U14 ( .A1(n944), .A2(n943), .A3(n942), .A4(n941), .ZN(N4481) );
  nd04d0 U15 ( .A1(n904), .A2(n903), .A3(n902), .A4(n901), .ZN(N4471) );
  nd04d0 U16 ( .A1(n744), .A2(n743), .A3(n742), .A4(n741), .ZN(N4494) );
  nd04d0 U17 ( .A1(n964), .A2(n963), .A3(n962), .A4(n961), .ZN(N4463) );
  nd04d0 U18 ( .A1(n882), .A2(n881), .A3(n880), .A4(n879), .ZN(N4483) );
  nd04d0 U19 ( .A1(n809), .A2(n808), .A3(n807), .A4(n806), .ZN(N4478) );
  nd04d0 U20 ( .A1(n721), .A2(n720), .A3(n719), .A4(n718), .ZN(
        mgmtsoc_ibus_ibus_dat_r[2]) );
  nd04d0 U21 ( .A1(n4683), .A2(n2476), .A3(n2475), .A4(n2474), .ZN(n2478) );
  nd04d0 U22 ( .A1(n459), .A2(n458), .A3(n457), .A4(n456), .ZN(n469) );
  nd04d0 U23 ( .A1(n5099), .A2(n5056), .A3(n5054), .A4(n5051), .ZN(n5057) );
  nd04d0 U24 ( .A1(mprj_adr_o[28]), .A2(n5716), .A3(n682), .A4(n681), .ZN(
        n1545) );
  nd04d0 U25 ( .A1(n1572), .A2(n1571), .A3(n1570), .A4(n1569), .ZN(n1582) );
  nd04d0 U26 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(n5049) );
  nd04d0 U27 ( .A1(n329), .A2(n328), .A3(mprj_adr_o[26]), .A4(mprj_adr_o[25]), 
        .ZN(n683) );
  nd04d0 U28 ( .A1(n1564), .A2(n1563), .A3(n1562), .A4(n1561), .ZN(n1583) );
  nd04d0 U29 ( .A1(n682), .A2(n5690), .A3(n5694), .A4(n346), .ZN(n352) );
  nd04d0 U30 ( .A1(n350), .A2(n5716), .A3(n5712), .A4(n367), .ZN(n351) );
  nd04d0 U31 ( .A1(n2793), .A2(n2792), .A3(n2791), .A4(n2790), .ZN(n2808) );
  nd04d0 U32 ( .A1(n2805), .A2(n2804), .A3(n2803), .A4(n2802), .ZN(n2807) );
  nd04d0 U33 ( .A1(n2763), .A2(n2762), .A3(n2761), .A4(n2760), .ZN(n2764) );
  nd04d0 U34 ( .A1(n2771), .A2(n2770), .A3(n2769), .A4(n2768), .ZN(n2777) );
  nd04d0 U35 ( .A1(n2786), .A2(n2785), .A3(n2784), .A4(n2783), .ZN(n2787) );
  nd04d0 U36 ( .A1(n2782), .A2(n2781), .A3(n2780), .A4(n2779), .ZN(n2788) );
  nd04d0 U37 ( .A1(n2775), .A2(n2774), .A3(n2773), .A4(n2772), .ZN(n2776) );
  nd04d0 U38 ( .A1(n2689), .A2(n2688), .A3(n2687), .A4(n2686), .ZN(n2690) );
  nd04d0 U39 ( .A1(n1898), .A2(n4881), .A3(n1897), .A4(n1896), .ZN(n1899) );
  nd04d0 U40 ( .A1(n1880), .A2(n1879), .A3(n1878), .A4(n1877), .ZN(n1881) );
  nd04d0 U41 ( .A1(n5108), .A2(n5107), .A3(n5106), .A4(n5105), .ZN(n5109) );
  nd04d0 U42 ( .A1(n5104), .A2(n5103), .A3(n5102), .A4(n5101), .ZN(n5110) );
  nd04d0 U43 ( .A1(n535), .A2(n534), .A3(n533), .A4(n532), .ZN(n1613) );
  nd04d0 U44 ( .A1(n2957), .A2(n2956), .A3(n2955), .A4(n2954), .ZN(n2965) );
  nd04d0 U45 ( .A1(n3017), .A2(n3016), .A3(n3015), .A4(n3014), .ZN(n3018) );
  nd04d0 U46 ( .A1(n3029), .A2(n3028), .A3(n3027), .A4(n3026), .ZN(n3044) );
  nd04d0 U47 ( .A1(n2939), .A2(n2938), .A3(n2937), .A4(n2936), .ZN(n2940) );
  nd04d0 U48 ( .A1(n358), .A2(n357), .A3(n1625), .A4(n356), .ZN(n1660) );
  nd04d0 U49 ( .A1(n2979), .A2(n2978), .A3(n2977), .A4(n2976), .ZN(n2980) );
  nd04d0 U50 ( .A1(n2989), .A2(n2988), .A3(n2987), .A4(n2986), .ZN(n2995) );
  nd04d0 U51 ( .A1(n2950), .A2(n2949), .A3(n2948), .A4(n2947), .ZN(n2951) );
  nd04d0 U52 ( .A1(n5301), .A2(n4640), .A3(n4641), .A4(n4642), .ZN(n4617) );
  nd04d0 U53 ( .A1(n2935), .A2(n2934), .A3(n2933), .A4(n2932), .ZN(n2941) );
  nd04d0 U54 ( .A1(n5949), .A2(n4765), .A3(n1249), .A4(n4768), .ZN(n1866) );
  nd04d0 U55 ( .A1(n5913), .A2(n4765), .A3(n5928), .A4(n1251), .ZN(n1867) );
  nd04d0 U56 ( .A1(n5932), .A2(n4765), .A3(n1249), .A4(n4769), .ZN(n1870) );
  nd04d0 U57 ( .A1(n304), .A2(n303), .A3(n302), .A4(n301), .ZN(n305) );
  nd04d0 U58 ( .A1(n404), .A2(n403), .A3(n402), .A4(n401), .ZN(n406) );
  nd02d0 U59 ( .A1(n613), .A2(n5912), .ZN(n541) );
  nr04d0 U60 ( .A1(mprj_adr_o[27]), .A2(mprj_adr_o[24]), .A3(mprj_adr_o[20]), 
        .A4(mprj_adr_o[21]), .ZN(n346) );
  nd03d0 U61 ( .A1(n613), .A2(n612), .A3(n5777), .ZN(n614) );
  nd02d0 U62 ( .A1(n5784), .A2(n661), .ZN(n5786) );
  nd03d0 U63 ( .A1(n2915), .A2(n2914), .A3(n2913), .ZN(n2930) );
  nd02d0 U64 ( .A1(n1903), .A2(n2373), .ZN(n729) );
  nr02d0 U65 ( .A1(n724), .A2(n2372), .ZN(n722) );
  nr02d0 U66 ( .A1(n1786), .A2(n729), .ZN(n824) );
  nd02d0 U67 ( .A1(n2474), .A2(n1829), .ZN(n2372) );
  nd02d0 U68 ( .A1(n1982), .A2(n2474), .ZN(n4960) );
  nr02d0 U69 ( .A1(n4811), .A2(n1783), .ZN(n2449) );
  nr02d0 U70 ( .A1(n1783), .A2(n4576), .ZN(n1805) );
  nd03d0 U71 ( .A1(n2614), .A2(n2620), .A3(n2613), .ZN(n2637) );
  nd03d0 U72 ( .A1(uart_tx_fifo_produce[3]), .A2(n2614), .A3(n2613), .ZN(n2608) );
  nd02d0 U73 ( .A1(n2621), .A2(n2620), .ZN(n2633) );
  nd02d0 U74 ( .A1(uart_tx_fifo_produce[3]), .A2(n2621), .ZN(n2605) );
  nd02d0 U75 ( .A1(uart_tx_fifo_produce[2]), .A2(n2615), .ZN(n2624) );
  nd02d0 U76 ( .A1(uart_tx_fifo_produce[2]), .A2(n2559), .ZN(n2591) );
  nr04d0 U77 ( .A1(mprj_adr_o[16]), .A2(mprj_adr_o[17]), .A3(mprj_adr_o[18]), 
        .A4(mprj_adr_o[19]), .ZN(n350) );
  nr04d0 U78 ( .A1(n5730), .A2(n5722), .A3(n352), .A4(n746), .ZN(n390) );
  nr03d0 U79 ( .A1(mprj_adr_o[8]), .A2(mprj_adr_o[9]), .A3(mprj_adr_o[10]), 
        .ZN(n389) );
  nr02d0 U80 ( .A1(mprj_adr_o[26]), .A2(mprj_adr_o[25]), .ZN(n682) );
  nd03d0 U81 ( .A1(n5730), .A2(n5722), .A3(n327), .ZN(n680) );
  nd02d0 U82 ( .A1(n308), .A2(n307), .ZN(n979) );
  nd02d0 U83 ( .A1(n1515), .A2(n5488), .ZN(n1513) );
  nd02d0 U84 ( .A1(n1895), .A2(n979), .ZN(n1532) );
  nd02d0 U85 ( .A1(n5490), .A2(dbg_uart_rx_rx), .ZN(n1524) );
  nd02d0 U86 ( .A1(n377), .A2(n376), .ZN(n5241) );
  nd02d0 U87 ( .A1(n1516), .A2(n5489), .ZN(n5342) );
  nr03d0 U88 ( .A1(n5611), .A2(n1327), .A3(mprj_adr_o[3]), .ZN(n726) );
  nd02d0 U89 ( .A1(n1764), .A2(mprj_adr_o[4]), .ZN(n1786) );
  nd02d0 U90 ( .A1(n723), .A2(mprj_adr_o[4]), .ZN(n727) );
  nd02d0 U91 ( .A1(n726), .A2(mprj_adr_o[4]), .ZN(n725) );
  nr02d0 U92 ( .A1(n469), .A2(n468), .ZN(n1205) );
  nr02d0 U93 ( .A1(mprj_adr_o[31]), .A2(mprj_adr_o[30]), .ZN(n367) );
  an02d0 U94 ( .A1(n979), .A2(n1888), .Z(mgmtsoc_dbus_dbus_ack) );
  nr02d0 U95 ( .A1(n1783), .A2(n4960), .ZN(n1794) );
  nd02d0 U96 ( .A1(n5784), .A2(n5783), .ZN(n5877) );
  an03d0 U97 ( .A1(n922), .A2(n921), .A3(n920), .Z(n923) );
  nd02d0 U98 ( .A1(n5862), .A2(n572), .ZN(n5900) );
  nd02d0 U99 ( .A1(n5862), .A2(n626), .ZN(n5905) );
  nd02d0 U100 ( .A1(n5862), .A2(n646), .ZN(n5911) );
  ad01d0 U101 ( .A(n5932), .B(n5931), .CI(n5930), .CO(n5937), .S(n5933) );
  ad01d0 U102 ( .A(n5913), .B(n5912), .CI(n5920), .CO(n5930), .S(n5919) );
  nd02d0 U103 ( .A1(n2013), .A2(mprj_dat_o[4]), .ZN(n4866) );
  an03d0 U104 ( .A1(n930), .A2(n929), .A3(n928), .Z(n931) );
  nd02d0 U105 ( .A1(n2013), .A2(mprj_dat_o[5]), .ZN(n2640) );
  nd02d0 U106 ( .A1(n2013), .A2(mprj_dat_o[3]), .ZN(n2625) );
  nr02d0 U107 ( .A1(n3060), .A2(n2655), .ZN(n2557) );
  nr02d0 U108 ( .A1(n1762), .A2(n1807), .ZN(n4579) );
  nr02d0 U109 ( .A1(n2462), .A2(n1807), .ZN(n1821) );
  nd02d0 U110 ( .A1(n1838), .A2(n1843), .ZN(n1845) );
  nd02d0 U111 ( .A1(n1843), .A2(n4952), .ZN(n1844) );
  nd02d0 U112 ( .A1(n2476), .A2(n4806), .ZN(n4810) );
  nd02d0 U113 ( .A1(n1903), .A2(n4806), .ZN(n1840) );
  nd03d0 U114 ( .A1(n4822), .A2(n5956), .A3(n4842), .ZN(n4834) );
  nd02d0 U115 ( .A1(n4812), .A2(n5956), .ZN(n4821) );
  nr04d0 U116 ( .A1(n5621), .A2(n724), .A3(n2372), .A4(n1762), .ZN(n945) );
  nr02d0 U117 ( .A1(n725), .A2(n729), .ZN(n919) );
  nr02d0 U118 ( .A1(n728), .A2(n727), .ZN(n947) );
  nd02d0 U119 ( .A1(litespiphy_state[0]), .A2(litespiphy_state[1]), .ZN(n4684)
         );
  nd02d0 U120 ( .A1(n723), .A2(n1765), .ZN(n1846) );
  nd02d0 U121 ( .A1(n726), .A2(n1765), .ZN(n1847) );
  nd02d0 U122 ( .A1(n2457), .A2(n2449), .ZN(n4959) );
  nd02d0 U123 ( .A1(n1829), .A2(n2466), .ZN(n4860) );
  nr02d0 U124 ( .A1(n4957), .A2(n4860), .ZN(n4861) );
  nd02d0 U125 ( .A1(n5955), .A2(n4870), .ZN(n4871) );
  nr03d0 U126 ( .A1(n5653), .A2(mprj_adr_o[14]), .A3(mprj_adr_o[15]), .ZN(
        n1829) );
  nr03d0 U127 ( .A1(n5645), .A2(n5649), .A3(n1327), .ZN(n1325) );
  nr03d0 U128 ( .A1(n5649), .A2(mprj_adr_o[11]), .A3(n1327), .ZN(n2474) );
  nd02d0 U129 ( .A1(n4998), .A2(n1903), .ZN(n3060) );
  nd03d0 U130 ( .A1(n5653), .A2(n5657), .A3(n5661), .ZN(n2470) );
  nr04d0 U131 ( .A1(mgmtsoc_dbus_dbus_sel[3]), .A2(mgmtsoc_dbus_dbus_sel[1]), 
        .A3(mgmtsoc_dbus_dbus_sel[0]), .A4(mprj_sel_o[2]), .ZN(n348) );
  nr02d0 U132 ( .A1(mprj_adr_o[13]), .A2(n369), .ZN(n1982) );
  nd03d0 U133 ( .A1(n2476), .A2(n1325), .A3(n1328), .ZN(n1976) );
  nd02d0 U134 ( .A1(n5288), .A2(n1981), .ZN(n1980) );
  nd02d0 U135 ( .A1(n1982), .A2(n1325), .ZN(n2655) );
  nd02d0 U136 ( .A1(n1839), .A2(n2449), .ZN(n2654) );
  nd02d0 U137 ( .A1(n5617), .A2(n723), .ZN(n2454) );
  nd02d0 U138 ( .A1(n4952), .A2(n2449), .ZN(n2334) );
  nd02d0 U139 ( .A1(n5617), .A2(n1764), .ZN(n2451) );
  nd02d0 U140 ( .A1(n4683), .A2(n2295), .ZN(n2300) );
  nd02d0 U141 ( .A1(n4683), .A2(n2183), .ZN(n2186) );
  nd02d0 U142 ( .A1(n4998), .A2(n4997), .ZN(n5001) );
  nr02d0 U143 ( .A1(n4960), .A2(n392), .ZN(n4997) );
  nd03d0 U144 ( .A1(n1982), .A2(n5649), .A3(mprj_adr_o[11]), .ZN(n4576) );
  nd03d0 U145 ( .A1(n4683), .A2(n1903), .A3(n1902), .ZN(n4575) );
  nr02d0 U146 ( .A1(n4811), .A2(n4810), .ZN(n4812) );
  nr02d0 U147 ( .A1(n3059), .A2(n2470), .ZN(n4806) );
  or02d0 U148 ( .A1(n4773), .A2(n4957), .Z(n4795) );
  nd02d0 U149 ( .A1(n5288), .A2(n4805), .ZN(n4797) );
  nd02d0 U150 ( .A1(n2560), .A2(n2620), .ZN(n2611) );
  nr02d0 U151 ( .A1(n2615), .A2(n2558), .ZN(n2559) );
  nr02d0 U152 ( .A1(n2594), .A2(n2613), .ZN(n2621) );
  nd03d0 U153 ( .A1(n2580), .A2(n2590), .A3(n2561), .ZN(n2569) );
  nd02d0 U154 ( .A1(n2148), .A2(n4580), .ZN(n2166) );
  nd02d0 U155 ( .A1(n4683), .A2(n1985), .ZN(n1989) );
  nr02d0 U156 ( .A1(n4576), .A2(n2334), .ZN(n1886) );
  nd02d0 U157 ( .A1(n4683), .A2(N6326), .ZN(n4957) );
  nd02d0 U158 ( .A1(n350), .A2(n390), .ZN(n349) );
  nd12d0 U159 ( .A1(n1532), .A2(n1515), .ZN(n5341) );
  nd02d0 U160 ( .A1(uartwishbonebridge_state[2]), .A2(n5296), .ZN(n1891) );
  nd03d0 U161 ( .A1(n5240), .A2(n5301), .A3(n5241), .ZN(n5286) );
  nd02d0 U162 ( .A1(uart_tx_fifo_level0[4]), .A2(n2563), .ZN(n2556) );
  nr02d0 U163 ( .A1(mgmtsoc_dbus_dbus_sel[2]), .A2(n378), .ZN(n354) );
  nd02d0 U164 ( .A1(n1900), .A2(n1895), .ZN(n1890) );
  nd02d0 U165 ( .A1(mprj_adr_o[29]), .A2(mprj_adr_o[28]), .ZN(n746) );
  nd02d0 U166 ( .A1(n1389), .A2(n1388), .ZN(mgmtsoc_ibus_ibus_dat_r[5]) );
  nd03d0 U167 ( .A1(n640), .A2(n639), .A3(n638), .ZN(n3137) );
  nd03d0 U168 ( .A1(n658), .A2(n657), .A3(n656), .ZN(n3136) );
  nd03d0 U169 ( .A1(n567), .A2(n566), .A3(n565), .ZN(n3135) );
  nd03d0 U170 ( .A1(n4683), .A2(n2466), .A3(n2465), .ZN(n2468) );
  nd03d0 U171 ( .A1(n4683), .A2(n1982), .A3(n2466), .ZN(n1984) );
  nd03d0 U172 ( .A1(n1911), .A2(gpioin4_pending_r), .A3(n5956), .ZN(n1910) );
  nd03d0 U173 ( .A1(n1943), .A2(csrbank17_edge0_w), .A3(n5956), .ZN(n1942) );
  nd03d0 U174 ( .A1(n4951), .A2(csrbank10_update_value0_w), .A3(n5956), .ZN(
        n4950) );
  nd03d0 U175 ( .A1(n4877), .A2(mgmtsoc_pending_r), .A3(n5301), .ZN(n4876) );
  nd03d0 U176 ( .A1(n2448), .A2(n6130), .A3(n5340), .ZN(n2447) );
  nr02d0 U177 ( .A1(n4957), .A2(n1826), .ZN(N5618) );
  an03d0 U178 ( .A1(n2013), .A2(hk_stb_o), .A3(N6304), .Z(N6326) );
  nr02d0 U179 ( .A1(n2516), .A2(n349), .ZN(N6304) );
  an02d0 U180 ( .A1(n1314), .A2(n1299), .Z(n4518) );
  an02d0 U181 ( .A1(n1314), .A2(n1302), .Z(n4519) );
  an02d0 U182 ( .A1(n1314), .A2(n1289), .Z(n4520) );
  an02d0 U183 ( .A1(n1314), .A2(n1287), .Z(n4521) );
  an02d0 U184 ( .A1(n1314), .A2(n1297), .Z(n4522) );
  an02d0 U185 ( .A1(n1314), .A2(n1310), .Z(n4524) );
  an02d0 U186 ( .A1(n1314), .A2(n1307), .Z(n4525) );
  an02d0 U187 ( .A1(n1314), .A2(n1312), .Z(n4527) );
  an02d0 U188 ( .A1(n1314), .A2(n1294), .Z(n4528) );
  an02d0 U189 ( .A1(n1314), .A2(n1291), .Z(n4529) );
  an02d0 U190 ( .A1(n1314), .A2(n1305), .Z(n4530) );
  an02d0 U191 ( .A1(n1314), .A2(n1285), .Z(n4532) );
  an02d0 U192 ( .A1(n5987), .A2(n1282), .Z(N5045) );
  an02d0 U193 ( .A1(n5987), .A2(n1273), .Z(N5044) );
  an02d0 U194 ( .A1(n5987), .A2(n1268), .Z(N5043) );
  an02d0 U195 ( .A1(n5987), .A2(n1246), .Z(N5042) );
  an02d0 U196 ( .A1(n5987), .A2(n1242), .Z(N5041) );
  an02d0 U197 ( .A1(n5987), .A2(n1235), .Z(N5040) );
  an02d0 U198 ( .A1(n5987), .A2(n1183), .Z(N5038) );
  an02d0 U199 ( .A1(n5987), .A2(n1145), .Z(N5033) );
  an02d0 U200 ( .A1(n5987), .A2(n1134), .Z(N5032) );
  an02d0 U201 ( .A1(n5987), .A2(n1117), .Z(N5030) );
  an02d0 U202 ( .A1(n5987), .A2(n1123), .Z(N5024) );
  an02d0 U203 ( .A1(n5987), .A2(n1125), .Z(N5023) );
  an02d0 U204 ( .A1(n5987), .A2(n1115), .Z(N5020) );
  an02d0 U205 ( .A1(n5987), .A2(n1113), .Z(N5019) );
  an02d0 U206 ( .A1(n5987), .A2(n1119), .Z(N5018) );
  an02d0 U207 ( .A1(n5987), .A2(n1121), .Z(N5017) );
  an02d0 U208 ( .A1(n5987), .A2(n1280), .Z(N5756) );
  aoi22d1 U209 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[2]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[2]), .ZN(n300) );
  nr03d0 U210 ( .A1(n5050), .A2(n746), .A3(n745), .ZN(mprj_cyc_o) );
  aoi22d1 U211 ( .A1(n3057), .A2(n3052), .B1(n3051), .B2(n3054), .ZN(n3725) );
  nd02d1 U212 ( .A1(n5955), .A2(n4581), .ZN(n4604) );
  inv0d2 U213 ( .I(n5492), .ZN(n5955) );
  inv0d2 U214 ( .I(uart_phy_rx_data[2]), .ZN(n3049) );
  inv0d2 U215 ( .I(n1890), .ZN(n342) );
  oai21d2 U216 ( .B1(n393), .B2(n5527), .A(n300), .ZN(mprj_adr_o[4]) );
  inv0d1 U217 ( .I(n661), .ZN(n659) );
  inv0d1 U218 ( .I(n5425), .ZN(n1451) );
  inv0d1 U219 ( .I(n4620), .ZN(n4566) );
  inv0d1 U220 ( .I(n2462), .ZN(n4998) );
  inv0d2 U221 ( .I(n4582), .ZN(n4808) );
  inv0d2 U222 ( .I(uart_phy_rx_data[7]), .ZN(n3055) );
  inv0d2 U223 ( .I(uart_phy_rx_data[5]), .ZN(n3052) );
  inv0d2 U224 ( .I(uart_phy_rx_data[3]), .ZN(n3050) );
  inv0d2 U225 ( .I(uart_phy_rx_data[1]), .ZN(n3048) );
  aoi21d4 U226 ( .B1(n5931), .B2(n541), .A(n545), .ZN(n5862) );
  nr02d2 U227 ( .A1(n5100), .A2(n1205), .ZN(n4678) );
  inv0d2 U228 ( .I(state), .ZN(n2022) );
  nd02d1 U229 ( .A1(n5340), .A2(n5327), .ZN(n5467) );
  buffd1 U230 ( .I(n6130), .Z(gpio_out_pad) );
  nr03d2 U231 ( .A1(n2616), .A2(n2615), .A3(n2608), .ZN(n2596) );
  nr03d2 U232 ( .A1(n979), .A2(n2516), .A3(n5050), .ZN(n1314) );
  inv0d1 U233 ( .I(litespi_tx_mux_sel), .ZN(n4685) );
  inv0d1 U234 ( .I(grant[1]), .ZN(n1900) );
  nr04d0 U235 ( .A1(mgmtsoc_litespimmap_burst_adr[28]), .A2(
        mgmtsoc_litespimmap_burst_adr[29]), .A3(n1560), .A4(n1559), .ZN(n1561)
         );
  nd04d0 U236 ( .A1(n1580), .A2(n1579), .A3(n1578), .A4(n1577), .ZN(n1581) );
  nr04d0 U237 ( .A1(n5172), .A2(n5168), .A3(n5164), .A4(n5160), .ZN(n5103) );
  nr04d0 U238 ( .A1(interface0_bank_bus_dat_r[1]), .A2(
        interface3_bank_bus_dat_r[1]), .A3(interface4_bank_bus_dat_r[1]), .A4(
        interface6_bank_bus_dat_r[1]), .ZN(n706) );
  nr03d0 U239 ( .A1(interface3_bank_bus_dat_r[3]), .A2(
        interface6_bank_bus_dat_r[3]), .A3(interface4_bank_bus_dat_r[3]), .ZN(
        n5346) );
  nr03d0 U240 ( .A1(interface3_bank_bus_dat_r[7]), .A2(
        interface6_bank_bus_dat_r[7]), .A3(interface4_bank_bus_dat_r[7]), .ZN(
        n5365) );
  nr04d0 U241 ( .A1(interface6_bank_bus_dat_r[10]), .A2(
        interface3_bank_bus_dat_r[10]), .A3(interface10_bank_bus_dat_r[10]), 
        .A4(interface9_bank_bus_dat_r[10]), .ZN(n5393) );
  nr04d0 U242 ( .A1(interface6_bank_bus_dat_r[14]), .A2(
        interface3_bank_bus_dat_r[14]), .A3(interface10_bank_bus_dat_r[14]), 
        .A4(interface9_bank_bus_dat_r[14]), .ZN(n5428) );
  nr04d0 U243 ( .A1(interface0_bank_bus_dat_r[19]), .A2(
        interface3_bank_bus_dat_r[19]), .A3(interface6_bank_bus_dat_r[19]), 
        .A4(interface10_bank_bus_dat_r[19]), .ZN(n1442) );
  nr04d0 U244 ( .A1(interface0_bank_bus_dat_r[24]), .A2(
        interface3_bank_bus_dat_r[24]), .A3(interface6_bank_bus_dat_r[24]), 
        .A4(interface10_bank_bus_dat_r[24]), .ZN(n1430) );
  nr04d0 U245 ( .A1(interface0_bank_bus_dat_r[29]), .A2(
        interface3_bank_bus_dat_r[29]), .A3(interface6_bank_bus_dat_r[29]), 
        .A4(interface10_bank_bus_dat_r[29]), .ZN(n1379) );
  nd12d0 U246 ( .A1(mgmtsoc_value[28]), .A2(n1699), .ZN(n1704) );
  nd12d0 U247 ( .A1(mgmtsoc_value[26]), .A2(n1693), .ZN(n1696) );
  nd12d0 U248 ( .A1(mgmtsoc_value[22]), .A2(n1681), .ZN(n1684) );
  nd12d0 U249 ( .A1(mgmtsoc_value[14]), .A2(n1656), .ZN(n1657) );
  nd12d0 U250 ( .A1(mgmtsoc_value[4]), .A2(n1625), .ZN(n1628) );
  nd04d0 U251 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(n363) );
  nr04d0 U252 ( .A1(n724), .A2(mprj_adr_o[5]), .A3(n2372), .A4(n1762), .ZN(
        n737) );
  nd04d0 U253 ( .A1(n515), .A2(n514), .A3(n513), .A4(n512), .ZN(n524) );
  nd12d0 U254 ( .A1(uart_phy_tx_phase[19]), .A2(n1476), .ZN(n1478) );
  nr02d0 U255 ( .A1(n5986), .A2(n1535), .ZN(n1522) );
  nd12d0 U256 ( .A1(dbg_uart_count[8]), .A2(n1088), .ZN(n2493) );
  nr02d0 U257 ( .A1(n1891), .A2(n1900), .ZN(n1515) );
  nd12d0 U258 ( .A1(dbg_uart_rx_phase[13]), .A2(n1070), .ZN(n1072) );
  nr02d0 U259 ( .A1(mprj_adr_o[9]), .A2(n525), .ZN(\RAM256/SEL0[0] ) );
  nr02d0 U260 ( .A1(n383), .A2(n382), .ZN(dff_we[0]) );
  nr02d0 U261 ( .A1(n4685), .A2(n4768), .ZN(n5932) );
  nr02d0 U262 ( .A1(n5938), .A2(n540), .ZN(n564) );
  nr02d0 U263 ( .A1(n2372), .A2(n1846), .ZN(n832) );
  nr02d0 U264 ( .A1(n2372), .A2(n1847), .ZN(n875) );
  nr02d0 U265 ( .A1(n5931), .A2(n541), .ZN(n545) );
  nd12d0 U266 ( .A1(n540), .A2(n5938), .ZN(n5778) );
  nd04d0 U267 ( .A1(n3041), .A2(n3040), .A3(n3039), .A4(n3038), .ZN(n3043) );
  nd04d0 U268 ( .A1(n2993), .A2(n2992), .A3(n2991), .A4(n2990), .ZN(n2994) );
  nd04d0 U269 ( .A1(n2963), .A2(n2962), .A3(n2961), .A4(n2960), .ZN(n2964) );
  nd04d0 U270 ( .A1(n2946), .A2(n2945), .A3(n2944), .A4(n2943), .ZN(n2952) );
  nr02d0 U271 ( .A1(n2451), .A2(n1807), .ZN(n1822) );
  nr02d0 U272 ( .A1(n1595), .A2(n4840), .ZN(n1598) );
  nr04d0 U273 ( .A1(n5922), .A2(n5913), .A3(n5932), .A4(n5949), .ZN(n5736) );
  nd03d0 U274 ( .A1(n1870), .A2(n1867), .A3(n1866), .ZN(n5735) );
  nr02d0 U275 ( .A1(n1660), .A2(n363), .ZN(n1614) );
  nr03d0 U276 ( .A1(n5951), .A2(n1262), .A3(n1261), .ZN(n5950) );
  nr02d0 U277 ( .A1(n2462), .A2(n729), .ZN(n937) );
  nr03d0 U278 ( .A1(n5614), .A2(mprj_adr_o[2]), .A3(n1327), .ZN(n723) );
  nd03d0 U279 ( .A1(n377), .A2(n5661), .A3(mprj_adr_o[14]), .ZN(n369) );
  nr02d0 U280 ( .A1(n5100), .A2(n4551), .ZN(n4620) );
  nr02d0 U281 ( .A1(n2584), .A2(n2583), .ZN(n2586) );
  nr02d0 U282 ( .A1(mprj_adr_o[10]), .A2(n353), .ZN(n355) );
  nd12d0 U283 ( .A1(count[4]), .A2(n1286), .ZN(n1296) );
  nd12d0 U284 ( .A1(count[6]), .A2(n701), .ZN(n1309) );
  nr02d0 U285 ( .A1(n1524), .A2(n1514), .ZN(n1529) );
  nd12d0 U286 ( .A1(dbg_uart_count[4]), .A2(n1100), .ZN(n1083) );
  nd12d0 U287 ( .A1(dbg_uart_count[12]), .A2(n1135), .ZN(n1168) );
  nr02d0 U288 ( .A1(dbg_uart_tx_phase[20]), .A2(n1751), .ZN(n1748) );
  nr02d0 U289 ( .A1(dbg_uart_tx_phase[7]), .A2(n1722), .ZN(n1725) );
  nr02d0 U290 ( .A1(n5050), .A2(n5049), .ZN(n5051) );
  nr02d0 U291 ( .A1(n5637), .A2(n709), .ZN(n5380) );
  nd04d0 U292 ( .A1(n1344), .A2(n1343), .A3(n1342), .A4(n1341), .ZN(n1345) );
  nr03d0 U293 ( .A1(n3011), .A2(n3010), .A3(n3009), .ZN(n3023) );
  nr04d0 U294 ( .A1(n2759), .A2(n2758), .A3(n2757), .A4(n2756), .ZN(n2766) );
  nr03d0 U295 ( .A1(n2975), .A2(n2974), .A3(n2973), .ZN(n2982) );
  nd12d0 U296 ( .A1(n5004), .A2(n5340), .ZN(n2298) );
  nr04d0 U297 ( .A1(n2842), .A2(n2841), .A3(n2840), .A4(n2839), .ZN(n2843) );
  nd12d0 U298 ( .A1(n4682), .A2(n4622), .ZN(n4660) );
  nr02d0 U299 ( .A1(n3085), .A2(n3089), .ZN(n4677) );
  nr03d0 U300 ( .A1(n5732), .A2(n4859), .A3(n4878), .ZN(n993) );
  nd03d0 U301 ( .A1(n1605), .A2(n1604), .A3(n1603), .ZN(n1609) );
  nd03d0 U302 ( .A1(n5649), .A2(n2465), .A3(mprj_adr_o[11]), .ZN(n1973) );
  nr02d0 U303 ( .A1(n1966), .A2(n4959), .ZN(n1968) );
  nr02d0 U304 ( .A1(n1952), .A2(n4959), .ZN(n1954) );
  nr02d0 U305 ( .A1(n1937), .A2(n4959), .ZN(n1939) );
  nd03d0 U306 ( .A1(n377), .A2(n5649), .A3(mprj_adr_o[11]), .ZN(n2469) );
  nr04d0 U307 ( .A1(n1327), .A2(n3060), .A3(mprj_adr_o[11]), .A4(
        mprj_adr_o[12]), .ZN(n2466) );
  nr02d0 U308 ( .A1(n1973), .A2(n2334), .ZN(n1972) );
  nr02d0 U309 ( .A1(n2451), .A2(n2461), .ZN(n2453) );
  nr02d0 U310 ( .A1(n4576), .A2(n4575), .ZN(n4578) );
  nd03d0 U311 ( .A1(n4574), .A2(n4572), .A3(n4607), .ZN(n4573) );
  nr03d0 U312 ( .A1(n2685), .A2(n2684), .A3(n2683), .ZN(n2692) );
  nr02d0 U313 ( .A1(n2669), .A2(n2668), .ZN(n2673) );
  nd04d0 U314 ( .A1(request[1]), .A2(n5340), .A3(n1893), .A4(n1901), .ZN(n1894) );
  nd12d0 U315 ( .A1(n406), .A2(n405), .ZN(n2497) );
  nr02d0 U316 ( .A1(n5100), .A2(n2874), .ZN(n1163) );
  nd04d0 U317 ( .A1(n713), .A2(n712), .A3(n711), .A4(n710), .ZN(
        mgmtsoc_ibus_ibus_dat_r[1]) );
  nd04d0 U318 ( .A1(n781), .A2(n780), .A3(n779), .A4(n778), .ZN(N4493) );
  nd04d0 U319 ( .A1(n954), .A2(n953), .A3(n952), .A4(n951), .ZN(N4492) );
  nd04d0 U320 ( .A1(n697), .A2(n696), .A3(n695), .A4(n694), .ZN(n3155) );
  nd04d0 U321 ( .A1(n978), .A2(n977), .A3(n976), .A4(n975), .ZN(N4491) );
  nd04d0 U322 ( .A1(n846), .A2(n845), .A3(n844), .A4(n843), .ZN(N4490) );
  nd04d0 U323 ( .A1(n874), .A2(n873), .A3(n872), .A4(n871), .ZN(N4489) );
  nd04d0 U324 ( .A1(n753), .A2(n752), .A3(n751), .A4(n750), .ZN(N4488) );
  nd03d0 U325 ( .A1(n561), .A2(n560), .A3(n559), .ZN(n3150) );
  nd03d0 U326 ( .A1(n632), .A2(n631), .A3(n630), .ZN(n3149) );
  nd04d0 U327 ( .A1(n839), .A2(n838), .A3(n837), .A4(n836), .ZN(N4485) );
  nd03d0 U328 ( .A1(n653), .A2(n652), .A3(n651), .ZN(n3148) );
  nd03d0 U329 ( .A1(n554), .A2(n553), .A3(n552), .ZN(n3147) );
  nd03d0 U330 ( .A1(n577), .A2(n576), .A3(n575), .ZN(n3146) );
  nd04d0 U331 ( .A1(n774), .A2(n773), .A3(n772), .A4(n771), .ZN(N4482) );
  nd03d0 U332 ( .A1(n620), .A2(n619), .A3(n618), .ZN(n3145) );
  nd03d0 U333 ( .A1(n603), .A2(n602), .A3(n601), .ZN(n3144) );
  nd03d0 U334 ( .A1(n589), .A2(n588), .A3(n587), .ZN(n3142) );
  nd03d0 U335 ( .A1(n636), .A2(n635), .A3(n634), .ZN(n3141) );
  nd04d0 U336 ( .A1(n897), .A2(n896), .A3(n895), .A4(n894), .ZN(N4477) );
  nd03d0 U337 ( .A1(n664), .A2(n663), .A3(n662), .ZN(n3140) );
  nd04d0 U338 ( .A1(n802), .A2(n801), .A3(n800), .A4(n799), .ZN(N4476) );
  nd03d0 U339 ( .A1(n581), .A2(n580), .A3(n579), .ZN(n3139) );
  nd04d0 U340 ( .A1(n926), .A2(n925), .A3(n924), .A4(n923), .ZN(N4475) );
  nd03d0 U341 ( .A1(n585), .A2(n584), .A3(n583), .ZN(n3138) );
  nr02d0 U342 ( .A1(n4867), .A2(n4860), .ZN(N4296) );
  nd04d0 U343 ( .A1(n823), .A2(n822), .A3(n821), .A4(n820), .ZN(N4467) );
  nd04d0 U344 ( .A1(n934), .A2(n933), .A3(n932), .A4(n931), .ZN(N4472) );
  nd04d0 U345 ( .A1(n816), .A2(n815), .A3(n814), .A4(n813), .ZN(N4468) );
  nr02d0 U346 ( .A1(n4865), .A2(n4860), .ZN(N4295) );
  nd04d0 U347 ( .A1(n853), .A2(n852), .A3(n851), .A4(n850), .ZN(N4466) );
  nd04d0 U348 ( .A1(n918), .A2(n917), .A3(n916), .A4(n915), .ZN(N4473) );
  nr02d0 U349 ( .A1(n4864), .A2(n4860), .ZN(N4294) );
  nd04d0 U350 ( .A1(n795), .A2(n794), .A3(n793), .A4(n792), .ZN(N4465) );
  nr02d0 U351 ( .A1(n1976), .A2(n1979), .ZN(N4997) );
  nr02d0 U352 ( .A1(n5100), .A2(n2662), .ZN(N5710) );
  nr02d0 U353 ( .A1(n1976), .A2(n1978), .ZN(N4996) );
  nd04d0 U354 ( .A1(n860), .A2(n859), .A3(n858), .A4(n857), .ZN(N4464) );
  nr02d0 U355 ( .A1(n4723), .A2(n4715), .ZN(N4271) );
  nr02d0 U356 ( .A1(n4723), .A2(n4716), .ZN(N4272) );
  nd04d0 U357 ( .A1(n911), .A2(n910), .A3(n909), .A4(n908), .ZN(N4469) );
  nd04d0 U358 ( .A1(n867), .A2(n866), .A3(n865), .A4(n864), .ZN(N4470) );
  nd04d0 U359 ( .A1(n767), .A2(n766), .A3(n765), .A4(n764), .ZN(N4474) );
  nr02d0 U360 ( .A1(n5100), .A2(n4880), .ZN(N5394) );
  nd04d0 U361 ( .A1(n788), .A2(n787), .A3(n786), .A4(n785), .ZN(N4487) );
  nd04d0 U362 ( .A1(n736), .A2(n735), .A3(n734), .A4(n733), .ZN(N4479) );
  nr02d0 U363 ( .A1(n2516), .A2(n1949), .ZN(N6231) );
  nr02d0 U364 ( .A1(n2516), .A2(n1934), .ZN(N6247) );
  nr03d0 U365 ( .A1(n5492), .A2(n2655), .A3(n2654), .ZN(N5711) );
  nr02d0 U366 ( .A1(n5492), .A2(n4951), .ZN(N5358) );
  nr02d0 U367 ( .A1(n1611), .A2(n4661), .ZN(n3663) );
  nr02d0 U368 ( .A1(n4957), .A2(n1848), .ZN(N5168) );
  nr02d0 U369 ( .A1(n2516), .A2(n672), .ZN(N6244) );
  inv0d0 U402 ( .I(grant[1]), .ZN(n393) );
  inv0d0 U403 ( .I(dbg_uart_wishbone_adr[2]), .ZN(n5527) );
  inv0d0 U404 ( .I(n393), .ZN(n341) );
  inv0d0 U405 ( .I(grant[0]), .ZN(n1895) );
  nr02d1 U406 ( .A1(n341), .A2(n1895), .ZN(n395) );
  inv0d0 U407 ( .I(n395), .ZN(n378) );
  inv0d2 U408 ( .I(n378), .ZN(n394) );
  nr04d0 U409 ( .A1(state), .A2(dff_bus_ack), .A3(dff2_bus_ack), .A4(
        mprj_ack_i), .ZN(n308) );
  nr02d0 U410 ( .A1(litespi_state[2]), .A2(litespi_state[1]), .ZN(n4845) );
  nd13d1 U411 ( .A1(litespi_state[0]), .A2(n4845), .A3(litespi_state[3]), .ZN(
        n1546) );
  nr03d0 U412 ( .A1(litespi_tx_mux_sel), .A2(n4684), .A3(n1546), .ZN(n5726) );
  buffd1 U413 ( .I(n5726), .Z(n5664) );
  or02d0 U414 ( .A1(count[14]), .A2(count[16]), .Z(n306) );
  nr04d0 U415 ( .A1(count[17]), .A2(count[19]), .A3(count[18]), .A4(count[2]), 
        .ZN(n304) );
  nr04d0 U416 ( .A1(count[9]), .A2(count[4]), .A3(count[5]), .A4(count[0]), 
        .ZN(n303) );
  nr04d0 U417 ( .A1(count[10]), .A2(count[8]), .A3(count[12]), .A4(count[3]), 
        .ZN(n302) );
  nr04d0 U418 ( .A1(count[11]), .A2(count[6]), .A3(count[7]), .A4(count[1]), 
        .ZN(n301) );
  or04d1 U419 ( .A1(count[15]), .A2(count[13]), .A3(n306), .A4(n305), .Z(n5425) );
  nr04d0 U420 ( .A1(n5664), .A2(n1451), .A3(hk_ack_i), .A4(
        mgmtsoc_vexriscv_debug_bus_ack), .ZN(n307) );
  nr02d0 U421 ( .A1(n341), .A2(n1532), .ZN(mgmtsoc_ibus_ibus_ack) );
  inv0d2 U422 ( .I(n378), .ZN(n1888) );
  aoi22d1 U423 ( .A1(n1888), .A2(mgmtsoc_dbus_dbus_adr[9]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[9]), .ZN(n309) );
  oaim21d1 U424 ( .B1(n341), .B2(dbg_uart_wishbone_adr[9]), .A(n309), .ZN(
        mprj_adr_o[11]) );
  inv0d0 U425 ( .I(dbg_uart_wishbone_adr[12]), .ZN(n5534) );
  aoi22d1 U426 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[12]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[12]), .ZN(n310) );
  oai21d1 U427 ( .B1(n1900), .B2(n5534), .A(n310), .ZN(mprj_adr_o[14]) );
  inv0d1 U428 ( .I(n393), .ZN(n397) );
  aoi22d1 U429 ( .A1(n397), .A2(dbg_uart_wishbone_adr[3]), .B1(n1888), .B2(
        mgmtsoc_dbus_dbus_adr[3]), .ZN(n311) );
  oai21d2 U430 ( .B1(mgmtsoc_ibus_ibus_adr[3]), .B2(n1890), .A(n311), .ZN(
        mprj_adr_o[5]) );
  inv0d0 U431 ( .I(request[0]), .ZN(n1893) );
  inv0d0 U432 ( .I(uartwishbonebridge_state[1]), .ZN(n5296) );
  aoi21d1 U433 ( .B1(n394), .B2(request[1]), .A(n1515), .ZN(n312) );
  oai21d1 U434 ( .B1(n1890), .B2(n1893), .A(n312), .ZN(hk_stb_o) );
  buffd1 U435 ( .I(rs232phy_rs232phyrx_state), .Z(n1200) );
  nd02d0 U436 ( .A1(n1200), .A2(uart_phy_rx_tick), .ZN(n3054) );
  inv0d0 U437 ( .I(n3054), .ZN(n3057) );
  nd02d0 U438 ( .A1(n3057), .A2(uart_phy_rx_count[0]), .ZN(n2889) );
  inv0d0 U439 ( .I(uart_phy_rx_count[3]), .ZN(n2890) );
  nr04d0 U440 ( .A1(uart_phy_rx_count[1]), .A2(uart_phy_rx_count[2]), .A3(
        n2889), .A4(n2890), .ZN(n2519) );
  inv0d0 U441 ( .I(uart_phy_rx_rx), .ZN(n3056) );
  buffd1 U442 ( .I(sys_rst), .Z(n4878) );
  buffd1 U443 ( .I(n4878), .Z(n5111) );
  inv0d2 U444 ( .I(n5111), .ZN(n5956) );
  aon211d1 U445 ( .C1(uart_phy_rx_rx_d), .C2(n3056), .B(n1200), .A(n4881), 
        .ZN(n313) );
  nr02d0 U446 ( .A1(n2519), .A2(n313), .ZN(n3869) );
  inv0d0 U447 ( .I(uartwishbonebridge_state[0]), .ZN(n5488) );
  oaim21d1 U448 ( .B1(n394), .B2(mgmtsoc_dbus_dbus_we), .A(n1513), .ZN(
        mprj_we_o) );
  inv0d0 U449 ( .I(dbg_uart_wishbone_adr[1]), .ZN(n5523) );
  aoi22d1 U450 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[1]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[1]), .ZN(n314) );
  oai21d1 U451 ( .B1(n393), .B2(n5523), .A(n314), .ZN(mprj_adr_o[3]) );
  aoi22d1 U452 ( .A1(n1888), .A2(mgmtsoc_dbus_dbus_adr[10]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[10]), .ZN(n315) );
  oaim21d1 U453 ( .B1(n341), .B2(dbg_uart_wishbone_adr[10]), .A(n315), .ZN(
        mprj_adr_o[12]) );
  inv0d0 U454 ( .I(dbg_uart_wishbone_adr[0]), .ZN(n5518) );
  aoi22d1 U455 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[0]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[0]), .ZN(n316) );
  oai21d1 U456 ( .B1(n1900), .B2(n5518), .A(n316), .ZN(mprj_adr_o[2]) );
  inv0d0 U457 ( .I(dbg_uart_wishbone_adr[20]), .ZN(n5600) );
  buffd1 U458 ( .I(n342), .Z(n344) );
  aoi22d1 U459 ( .A1(n1888), .A2(mgmtsoc_dbus_dbus_adr[20]), .B1(n344), .B2(
        mgmtsoc_ibus_ibus_adr[20]), .ZN(n317) );
  oai21d1 U460 ( .B1(n1900), .B2(n5600), .A(n317), .ZN(mprj_adr_o[22]) );
  aoi22d1 U461 ( .A1(n1888), .A2(mgmtsoc_dbus_dbus_adr[21]), .B1(n344), .B2(
        mgmtsoc_ibus_ibus_adr[21]), .ZN(n318) );
  oaim21d1 U462 ( .B1(n341), .B2(dbg_uart_wishbone_adr[21]), .A(n318), .ZN(
        mprj_adr_o[23]) );
  inv0d0 U463 ( .I(dbg_uart_wishbone_adr[27]), .ZN(n5594) );
  aoi22d1 U464 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[27]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[27]), .ZN(n319) );
  oai21d1 U465 ( .B1(n393), .B2(n5594), .A(n319), .ZN(mprj_adr_o[29]) );
  inv0d0 U466 ( .I(dbg_uart_wishbone_adr[26]), .ZN(n5589) );
  aoi22d1 U467 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[26]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[26]), .ZN(n320) );
  oai21d1 U468 ( .B1(n1900), .B2(n5589), .A(n320), .ZN(mprj_adr_o[28]) );
  inv0d0 U469 ( .I(dbg_uart_wishbone_adr[29]), .ZN(n5608) );
  aoi22d1 U470 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[29]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[29]), .ZN(n321) );
  oai21d1 U471 ( .B1(n1900), .B2(n5608), .A(n321), .ZN(mprj_adr_o[31]) );
  aoi22d1 U472 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[28]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[28]), .ZN(n322) );
  oaim21d1 U473 ( .B1(n341), .B2(dbg_uart_wishbone_adr[28]), .A(n322), .ZN(
        mprj_adr_o[30]) );
  inv0d0 U474 ( .I(dbg_uart_wishbone_adr[25]), .ZN(n5585) );
  aoi22d1 U475 ( .A1(n1888), .A2(mgmtsoc_dbus_dbus_adr[25]), .B1(n344), .B2(
        mgmtsoc_ibus_ibus_adr[25]), .ZN(n323) );
  oai21d1 U476 ( .B1(n1900), .B2(n5585), .A(n323), .ZN(mprj_adr_o[27]) );
  inv0d0 U477 ( .I(dbg_uart_wishbone_adr[22]), .ZN(n5573) );
  aoi22d1 U478 ( .A1(n1888), .A2(mgmtsoc_dbus_dbus_adr[22]), .B1(n344), .B2(
        mgmtsoc_ibus_ibus_adr[22]), .ZN(n324) );
  oai21d1 U479 ( .B1(n1900), .B2(n5573), .A(n324), .ZN(mprj_adr_o[24]) );
  inv0d0 U480 ( .I(dbg_uart_wishbone_adr[24]), .ZN(n5581) );
  aoi22d1 U481 ( .A1(n1888), .A2(mgmtsoc_dbus_dbus_adr[24]), .B1(n344), .B2(
        mgmtsoc_ibus_ibus_adr[24]), .ZN(n325) );
  oai21d1 U482 ( .B1(n1900), .B2(n5581), .A(n325), .ZN(mprj_adr_o[26]) );
  inv0d0 U483 ( .I(dbg_uart_wishbone_adr[23]), .ZN(n5577) );
  aoi22d1 U484 ( .A1(n1888), .A2(mgmtsoc_dbus_dbus_adr[23]), .B1(n344), .B2(
        mgmtsoc_ibus_ibus_adr[23]), .ZN(n326) );
  oai21d1 U485 ( .B1(n1900), .B2(n5577), .A(n326), .ZN(mprj_adr_o[25]) );
  inv0d0 U486 ( .I(hk_stb_o), .ZN(n5050) );
  nr02d0 U487 ( .A1(mprj_adr_o[22]), .A2(mprj_adr_o[23]), .ZN(n329) );
  inv0d0 U488 ( .I(mprj_adr_o[29]), .ZN(n5716) );
  inv0d0 U489 ( .I(mprj_adr_o[31]), .ZN(n5730) );
  inv0d0 U490 ( .I(mprj_adr_o[30]), .ZN(n5722) );
  nr02d0 U491 ( .A1(mprj_adr_o[27]), .A2(mprj_adr_o[24]), .ZN(n327) );
  nr03d0 U492 ( .A1(n5716), .A2(mprj_adr_o[28]), .A3(n680), .ZN(n328) );
  nr02d0 U493 ( .A1(n5050), .A2(n683), .ZN(hk_cyc_o) );
  aoi22d1 U494 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[14]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[14]), .ZN(n330) );
  oaim21d1 U495 ( .B1(n341), .B2(dbg_uart_wishbone_adr[14]), .A(n330), .ZN(
        mprj_adr_o[16]) );
  inv0d0 U496 ( .I(dbg_uart_wishbone_adr[15]), .ZN(n5545) );
  aoi22d1 U497 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[15]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[15]), .ZN(n331) );
  oai21d1 U498 ( .B1(n1900), .B2(n5545), .A(n331), .ZN(mprj_adr_o[17]) );
  inv0d0 U499 ( .I(dbg_uart_wishbone_adr[16]), .ZN(n5549) );
  aoi22d1 U500 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[16]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[16]), .ZN(n332) );
  oai21d1 U501 ( .B1(n393), .B2(n5549), .A(n332), .ZN(mprj_adr_o[18]) );
  inv0d0 U502 ( .I(dbg_uart_wishbone_adr[17]), .ZN(n5553) );
  aoi22d1 U503 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[17]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[17]), .ZN(n333) );
  oai21d1 U504 ( .B1(n393), .B2(n5553), .A(n333), .ZN(mprj_adr_o[19]) );
  inv0d0 U505 ( .I(dbg_uart_wishbone_adr[18]), .ZN(n5557) );
  aoi22d1 U506 ( .A1(n1888), .A2(mgmtsoc_dbus_dbus_adr[18]), .B1(n344), .B2(
        mgmtsoc_ibus_ibus_adr[18]), .ZN(n334) );
  oai21d1 U507 ( .B1(n1900), .B2(n5557), .A(n334), .ZN(mprj_adr_o[20]) );
  aoi22d1 U508 ( .A1(n1888), .A2(mgmtsoc_dbus_dbus_adr[19]), .B1(n344), .B2(
        mgmtsoc_ibus_ibus_adr[19]), .ZN(n335) );
  oaim21d1 U509 ( .B1(n341), .B2(dbg_uart_wishbone_adr[19]), .A(n335), .ZN(
        mprj_adr_o[21]) );
  aoi22d1 U510 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[5]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[5]), .ZN(n336) );
  oaim21d1 U511 ( .B1(n397), .B2(dbg_uart_wishbone_adr[5]), .A(n336), .ZN(
        mprj_adr_o[7]) );
  aoi22d1 U512 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[4]), .B1(n344), .B2(
        mgmtsoc_ibus_ibus_adr[4]), .ZN(n337) );
  oaim21d1 U513 ( .B1(n397), .B2(dbg_uart_wishbone_adr[4]), .A(n337), .ZN(
        mprj_adr_o[6]) );
  inv0d0 U514 ( .I(dbg_uart_wishbone_adr[6]), .ZN(n5541) );
  aoi22d1 U515 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[6]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[6]), .ZN(n338) );
  oai21d1 U516 ( .B1(n393), .B2(n5541), .A(n338), .ZN(mprj_adr_o[8]) );
  aoi22d1 U517 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[7]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[7]), .ZN(n339) );
  oaim21d1 U518 ( .B1(n397), .B2(dbg_uart_wishbone_adr[7]), .A(n339), .ZN(
        mprj_adr_o[9]) );
  aoi22d1 U519 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[8]), .B1(n344), .B2(
        mgmtsoc_ibus_ibus_adr[8]), .ZN(n340) );
  oaim21d1 U520 ( .B1(n341), .B2(dbg_uart_wishbone_adr[8]), .A(n340), .ZN(
        mprj_adr_o[10]) );
  inv0d0 U521 ( .I(dbg_uart_wishbone_adr[11]), .ZN(n5561) );
  aoi22d1 U522 ( .A1(n1888), .A2(mgmtsoc_dbus_dbus_adr[11]), .B1(n342), .B2(
        mgmtsoc_ibus_ibus_adr[11]), .ZN(n343) );
  oai21d1 U523 ( .B1(n1900), .B2(n5561), .A(n343), .ZN(mprj_adr_o[13]) );
  inv0d0 U524 ( .I(dbg_uart_wishbone_adr[13]), .ZN(n5568) );
  aoi22d1 U525 ( .A1(n394), .A2(mgmtsoc_dbus_dbus_adr[13]), .B1(n344), .B2(
        mgmtsoc_ibus_ibus_adr[13]), .ZN(n345) );
  oai21d1 U526 ( .B1(n1900), .B2(n5568), .A(n345), .ZN(mprj_adr_o[15]) );
  inv0d0 U527 ( .I(mprj_adr_o[2]), .ZN(n5611) );
  inv0d0 U528 ( .I(mprj_adr_o[3]), .ZN(n5614) );
  inv0d0 U529 ( .I(mprj_adr_o[4]), .ZN(n5617) );
  inv0d0 U530 ( .I(mprj_adr_o[22]), .ZN(n5690) );
  inv0d0 U531 ( .I(mprj_adr_o[23]), .ZN(n5694) );
  nr03d0 U532 ( .A1(state), .A2(n5050), .A3(n349), .ZN(n377) );
  inv0d0 U533 ( .I(n377), .ZN(n1327) );
  aoi31d1 U534 ( .B1(n5611), .B2(n5614), .B3(n5617), .A(n1327), .ZN(n2462) );
  inv0d0 U535 ( .I(mprj_adr_o[7]), .ZN(n5629) );
  inv0d0 U536 ( .I(mprj_adr_o[6]), .ZN(n5625) );
  aoi31d1 U537 ( .B1(n5629), .B2(n5625), .B3(n389), .A(n1327), .ZN(n724) );
  aoi21d1 U538 ( .B1(n377), .B2(mprj_adr_o[5]), .A(n724), .ZN(n1903) );
  inv0d0 U539 ( .I(mprj_adr_o[13]), .ZN(n5653) );
  inv0d0 U540 ( .I(mprj_adr_o[14]), .ZN(n5657) );
  inv0d0 U541 ( .I(mprj_adr_o[15]), .ZN(n5661) );
  inv0d0 U542 ( .I(mprj_adr_o[12]), .ZN(n5649) );
  inv0d0 U543 ( .I(debug_mode), .ZN(n347) );
  nr04d0 U544 ( .A1(n3060), .A2(n2470), .A3(n2469), .A4(n347), .ZN(N4141) );
  inv0d0 U545 ( .I(n354), .ZN(mprj_sel_o[2]) );
  buffd1 U546 ( .I(n4878), .Z(n5492) );
  inv0d0 U547 ( .I(mprj_adr_o[11]), .ZN(n5645) );
  nd03d0 U548 ( .A1(n5611), .A2(mprj_adr_o[4]), .A3(n5614), .ZN(n1762) );
  inv0d1 U549 ( .I(n1762), .ZN(n1839) );
  inv0d0 U550 ( .I(mprj_we_o), .ZN(n5097) );
  nr02d1 U551 ( .A1(n5097), .A2(n348), .ZN(n4683) );
  inv0d0 U552 ( .I(n4683), .ZN(n4811) );
  inv0d0 U553 ( .I(n1903), .ZN(n1783) );
  buffd1 U554 ( .I(n4878), .Z(n2516) );
  buffd1 U555 ( .I(n2022), .Z(n2013) );
  inv0d0 U556 ( .I(mprj_adr_o[10]), .ZN(n5641) );
  nr03d0 U557 ( .A1(mprj_adr_o[11]), .A2(mprj_adr_o[12]), .A3(n2470), .ZN(n388) );
  inv0d0 U558 ( .I(n388), .ZN(n376) );
  inv0d0 U559 ( .I(mprj_adr_o[28]), .ZN(n5712) );
  nr03d0 U560 ( .A1(n352), .A2(n376), .A3(n351), .ZN(n368) );
  nd02d0 U561 ( .A1(n368), .A2(hk_stb_o), .ZN(n353) );
  nr03d0 U562 ( .A1(n5641), .A2(mprj_adr_o[9]), .A3(n353), .ZN(dff2_en) );
  nd02d0 U563 ( .A1(dff2_en), .A2(mprj_we_o), .ZN(n381) );
  nr02d0 U564 ( .A1(n354), .A2(n381), .ZN(dff2_we[2]) );
  nd02d0 U565 ( .A1(n355), .A2(mprj_we_o), .ZN(n383) );
  nr02d0 U566 ( .A1(n354), .A2(n383), .ZN(dff_we[2]) );
  inv0d0 U567 ( .I(n355), .ZN(n525) );
  buffd1 U568 ( .I(n4878), .Z(n5100) );
  nr04d0 U569 ( .A1(mgmtsoc_value[11]), .A2(mgmtsoc_value[10]), .A3(
        mgmtsoc_value[9]), .A4(mgmtsoc_value[8]), .ZN(n358) );
  nr04d0 U570 ( .A1(mgmtsoc_value[15]), .A2(mgmtsoc_value[14]), .A3(
        mgmtsoc_value[13]), .A4(mgmtsoc_value[12]), .ZN(n357) );
  nr04d0 U571 ( .A1(mgmtsoc_value[3]), .A2(mgmtsoc_value[2]), .A3(
        mgmtsoc_value[1]), .A4(mgmtsoc_value[0]), .ZN(n1625) );
  nr04d0 U572 ( .A1(mgmtsoc_value[7]), .A2(mgmtsoc_value[6]), .A3(
        mgmtsoc_value[5]), .A4(mgmtsoc_value[4]), .ZN(n356) );
  nr04d0 U573 ( .A1(mgmtsoc_value[27]), .A2(mgmtsoc_value[26]), .A3(
        mgmtsoc_value[25]), .A4(mgmtsoc_value[24]), .ZN(n362) );
  nr04d0 U574 ( .A1(mgmtsoc_value[31]), .A2(mgmtsoc_value[30]), .A3(
        mgmtsoc_value[29]), .A4(mgmtsoc_value[28]), .ZN(n361) );
  nr04d0 U575 ( .A1(mgmtsoc_value[19]), .A2(mgmtsoc_value[18]), .A3(
        mgmtsoc_value[17]), .A4(mgmtsoc_value[16]), .ZN(n360) );
  nr04d0 U576 ( .A1(mgmtsoc_value[23]), .A2(mgmtsoc_value[22]), .A3(
        mgmtsoc_value[21]), .A4(mgmtsoc_value[20]), .ZN(n359) );
  inv0d0 U577 ( .I(n1614), .ZN(n4880) );
  nd02d0 U578 ( .A1(dbg_uart_rx_tick), .A2(dbg_uart_rx_count[0]), .ZN(n2872)
         );
  inv0d0 U579 ( .I(dbg_uart_rx_count[1]), .ZN(n364) );
  nr02d0 U580 ( .A1(n2872), .A2(n364), .ZN(n2873) );
  inv0d0 U581 ( .I(uartwishbonebridge_rs232phyrx_state), .ZN(n2874) );
  aoi211d1 U582 ( .C1(n2872), .C2(n364), .A(n2873), .B(n2874), .ZN(n3880) );
  inv0d0 U583 ( .I(n3880), .ZN(n365) );
  inv0d0 U584 ( .I(dbg_uart_rx_count[3]), .ZN(n2876) );
  nr04d0 U585 ( .A1(dbg_uart_rx_count[2]), .A2(n365), .A3(n2872), .A4(n2876), 
        .ZN(n5490) );
  inv0d0 U586 ( .I(dbg_uart_rx_rx), .ZN(n2879) );
  inv0d2 U587 ( .I(n5100), .ZN(n5319) );
  aon211d1 U588 ( .C1(dbg_uart_rx_rx_d), .C2(n2879), .B(
        uartwishbonebridge_rs232phyrx_state), .A(n5319), .ZN(n366) );
  nr02d0 U589 ( .A1(n5490), .A2(n366), .ZN(n3882) );
  inv0d0 U590 ( .I(n367), .ZN(n745) );
  nr03d0 U591 ( .A1(n5492), .A2(n746), .A3(n745), .ZN(N6302) );
  inv0d1 U592 ( .I(n5111), .ZN(n4881) );
  nd02d0 U593 ( .A1(n368), .A2(n5301), .ZN(n391) );
  nr03d0 U594 ( .A1(n5641), .A2(mprj_adr_o[9]), .A3(n391), .ZN(N6300) );
  nr02d0 U595 ( .A1(n5653), .A2(n369), .ZN(n2465) );
  nd02d0 U596 ( .A1(n1325), .A2(n2465), .ZN(n1959) );
  nr03d0 U597 ( .A1(n5492), .A2(n1959), .A3(n2654), .ZN(N6275) );
  inv0d1 U598 ( .I(n725), .ZN(n1902) );
  inv0d0 U599 ( .I(csrbank17_in_w), .ZN(n670) );
  inv0d0 U600 ( .I(csrbank17_mode0_w), .ZN(n1947) );
  aoi22d1 U601 ( .A1(csrbank17_mode0_w), .A2(gpioin4_gpioin4_in_pads_n_d), 
        .B1(csrbank17_edge0_w), .B2(n1947), .ZN(n370) );
  mx02d1 U602 ( .I0(csrbank17_in_w), .I1(n670), .S(n370), .Z(n1941) );
  nr02d0 U603 ( .A1(n5611), .A2(n5614), .ZN(n1764) );
  aoi22d1 U604 ( .A1(n4998), .A2(csrbank17_in_w), .B1(n1839), .B2(gpioin4_i01), 
        .ZN(n373) );
  inv0d0 U605 ( .I(n2454), .ZN(n4952) );
  inv0d0 U606 ( .I(n726), .ZN(n371) );
  nr02d1 U607 ( .A1(mprj_adr_o[4]), .A2(n371), .ZN(n2457) );
  aoi22d1 U608 ( .A1(n4952), .A2(csrbank17_edge0_w), .B1(csrbank17_mode0_w), 
        .B2(n2457), .ZN(n372) );
  oai211d1 U609 ( .C1(n1941), .C2(n2451), .A(n373), .B(n372), .ZN(n374) );
  nr03d0 U610 ( .A1(n5661), .A2(mprj_adr_o[14]), .A3(mprj_adr_o[13]), .ZN(
        n1328) );
  inv0d0 U611 ( .I(n1328), .ZN(n1326) );
  nr02d0 U612 ( .A1(n1326), .A2(n2469), .ZN(n1944) );
  aon211d1 U613 ( .C1(n1902), .C2(gpioin4_i02), .B(n374), .A(n1944), .ZN(n375)
         );
  nr02d0 U614 ( .A1(n1783), .A2(n375), .ZN(N4950) );
  inv0d0 U615 ( .I(n3060), .ZN(n2476) );
  nd02d0 U616 ( .A1(n2476), .A2(n5241), .ZN(n1848) );
  nr02d0 U617 ( .A1(n378), .A2(mgmtsoc_dbus_dbus_sel[0]), .ZN(n382) );
  inv0d0 U618 ( .I(n382), .ZN(mprj_sel_o[0]) );
  nr02d0 U619 ( .A1(n378), .A2(mgmtsoc_dbus_dbus_sel[3]), .ZN(n379) );
  inv0d0 U620 ( .I(n379), .ZN(mprj_sel_o[3]) );
  inv0d0 U621 ( .I(n2451), .ZN(n1838) );
  inv0d0 U622 ( .I(n1325), .ZN(n3059) );
  inv0d0 U623 ( .I(n1840), .ZN(n1843) );
  inv0d0 U624 ( .I(mgmtsoc_master_rxtx_w[24]), .ZN(n4711) );
  nr02d0 U625 ( .A1(n1845), .A2(n4711), .ZN(N4267) );
  inv0d0 U626 ( .I(n1805), .ZN(n1807) );
  inv0d0 U627 ( .I(n1821), .ZN(n1826) );
  nr02d0 U628 ( .A1(n378), .A2(mgmtsoc_dbus_dbus_sel[1]), .ZN(n380) );
  inv0d0 U629 ( .I(n380), .ZN(mprj_sel_o[1]) );
  aoi22d1 U630 ( .A1(n397), .A2(dbg_uart_wishbone_dat_w[2]), .B1(n1888), .B2(
        mgmtsoc_dbus_dbus_dat_w[2]), .ZN(n5060) );
  inv0d0 U631 ( .I(n5060), .ZN(mprj_dat_o[2]) );
  inv0d0 U632 ( .I(n393), .ZN(n396) );
  aoi22d1 U633 ( .A1(n396), .A2(dbg_uart_wishbone_dat_w[6]), .B1(n395), .B2(
        mgmtsoc_dbus_dbus_dat_w[6]), .ZN(n5064) );
  inv0d0 U634 ( .I(n5064), .ZN(mprj_dat_o[6]) );
  aoi22d1 U635 ( .A1(n397), .A2(dbg_uart_wishbone_dat_w[1]), .B1(n1888), .B2(
        mgmtsoc_dbus_dbus_dat_w[1]), .ZN(n5059) );
  inv0d0 U636 ( .I(n5059), .ZN(mprj_dat_o[1]) );
  aoi22d1 U637 ( .A1(n397), .A2(dbg_uart_wishbone_dat_w[3]), .B1(n1888), .B2(
        mgmtsoc_dbus_dbus_dat_w[3]), .ZN(n5061) );
  inv0d0 U638 ( .I(n5061), .ZN(mprj_dat_o[3]) );
  aoi22d1 U639 ( .A1(n397), .A2(dbg_uart_wishbone_dat_w[0]), .B1(n1888), .B2(
        mgmtsoc_dbus_dbus_dat_w[0]), .ZN(n5058) );
  inv0d0 U640 ( .I(n5058), .ZN(mprj_dat_o[0]) );
  aoi22d1 U641 ( .A1(n396), .A2(dbg_uart_wishbone_dat_w[7]), .B1(n1888), .B2(
        mgmtsoc_dbus_dbus_dat_w[7]), .ZN(n5065) );
  inv0d0 U642 ( .I(n5065), .ZN(mprj_dat_o[7]) );
  aoi22d1 U643 ( .A1(n396), .A2(dbg_uart_wishbone_dat_w[5]), .B1(n395), .B2(
        mgmtsoc_dbus_dbus_dat_w[5]), .ZN(n5063) );
  inv0d0 U644 ( .I(n5063), .ZN(mprj_dat_o[5]) );
  aoi22d1 U645 ( .A1(n397), .A2(dbg_uart_wishbone_dat_w[4]), .B1(n1888), .B2(
        mgmtsoc_dbus_dbus_dat_w[4]), .ZN(n5062) );
  inv0d0 U646 ( .I(n5062), .ZN(mprj_dat_o[4]) );
  nr02d0 U647 ( .A1(n379), .A2(n381), .ZN(dff2_we[3]) );
  nr02d0 U648 ( .A1(n379), .A2(n383), .ZN(dff_we[3]) );
  nr02d0 U649 ( .A1(n380), .A2(n381), .ZN(dff2_we[1]) );
  nr02d0 U650 ( .A1(n380), .A2(n383), .ZN(dff_we[1]) );
  nr02d0 U651 ( .A1(n382), .A2(n381), .ZN(dff2_we[0]) );
  inv0d0 U652 ( .I(mprj_adr_o[9]), .ZN(n5637) );
  nr02d0 U653 ( .A1(n5637), .A2(n525), .ZN(\RAM256/SEL0[1] ) );
  buffd1 U654 ( .I(core_clk), .Z(n6129) );
  buffd1 U655 ( .I(n6129), .Z(n6110) );
  buffd1 U656 ( .I(n6110), .Z(n6105) );
  buffd1 U657 ( .I(n6105), .Z(n6123) );
  buffd1 U658 ( .I(n6123), .Z(n6121) );
  buffd1 U659 ( .I(n6121), .Z(n6122) );
  buffd1 U660 ( .I(n6122), .Z(n6085) );
  buffd1 U661 ( .I(n6085), .Z(n6100) );
  buffd1 U662 ( .I(n6100), .Z(n6101) );
  buffd1 U663 ( .I(n6101), .Z(n6047) );
  buffd1 U664 ( .I(n6047), .Z(n6128) );
  buffd1 U665 ( .I(n6128), .Z(n6111) );
  nr02d0 U666 ( .A1(n5100), .A2(n3056), .ZN(N5704) );
  inv0d0 U667 ( .I(csrbank16_in_w), .ZN(n669) );
  nr02d0 U668 ( .A1(n5100), .A2(n669), .ZN(N6228) );
  inv0d0 U669 ( .I(\uart_status_status[1] ), .ZN(n2662) );
  inv0d0 U670 ( .I(uart_tx_fifo_level0[2]), .ZN(n2580) );
  inv0d0 U671 ( .I(uart_tx_fifo_level0[1]), .ZN(n2590) );
  inv0d0 U672 ( .I(uart_tx_fifo_level0[0]), .ZN(n2561) );
  nr02d0 U673 ( .A1(n2569), .A2(uart_tx_fifo_level0[3]), .ZN(n2563) );
  inv0d0 U674 ( .I(n2556), .ZN(n2664) );
  nr02d0 U675 ( .A1(n5100), .A2(n2664), .ZN(N5707) );
  nd02d0 U676 ( .A1(csrbank15_edge0_w), .A2(n4881), .ZN(n384) );
  nr02d0 U677 ( .A1(csrbank15_mode0_w), .A2(n384), .ZN(N6223) );
  inv0d1 U678 ( .I(n5492), .ZN(n5288) );
  nd02d0 U679 ( .A1(csrbank13_edge0_w), .A2(n5288), .ZN(n385) );
  nr02d0 U680 ( .A1(csrbank13_mode0_w), .A2(n385), .ZN(N6207) );
  nd02d0 U681 ( .A1(csrbank14_edge0_w), .A2(n5956), .ZN(n386) );
  nr02d0 U682 ( .A1(csrbank14_mode0_w), .A2(n386), .ZN(N6215) );
  inv0d0 U683 ( .I(mprj_adr_o[16]), .ZN(n5666) );
  inv0d0 U684 ( .I(mprj_adr_o[17]), .ZN(n5670) );
  inv0d0 U685 ( .I(mprj_adr_o[18]), .ZN(n5674) );
  inv0d0 U686 ( .I(mprj_adr_o[19]), .ZN(n5678) );
  nr04d0 U687 ( .A1(n5666), .A2(n5670), .A3(n5674), .A4(n5678), .ZN(n387) );
  nr02d0 U688 ( .A1(n2516), .A2(n5049), .ZN(N6298) );
  nr02d0 U689 ( .A1(mprj_adr_o[10]), .A2(n391), .ZN(N6299) );
  inv0d0 U690 ( .I(n727), .ZN(n1806) );
  inv0d0 U691 ( .I(n2449), .ZN(n392) );
  nd02d0 U692 ( .A1(n1806), .A2(n4997), .ZN(n4877) );
  nr02d0 U693 ( .A1(n5492), .A2(n4877), .ZN(N5395) );
  nr02d0 U694 ( .A1(n5100), .A2(n2879), .ZN(N5758) );
  nd02d0 U695 ( .A1(n1838), .A2(n4997), .ZN(n4951) );
  aoi22d1 U696 ( .A1(grant[1]), .A2(dbg_uart_wishbone_dat_w[22]), .B1(n395), 
        .B2(mgmtsoc_dbus_dbus_dat_w[22]), .ZN(n5081) );
  inv0d0 U697 ( .I(n5081), .ZN(mprj_dat_o[22]) );
  aoi22d1 U698 ( .A1(grant[1]), .A2(dbg_uart_wishbone_dat_w[26]), .B1(n394), 
        .B2(mgmtsoc_dbus_dbus_dat_w[26]), .ZN(n5086) );
  inv0d0 U699 ( .I(n5086), .ZN(mprj_dat_o[26]) );
  aoi22d1 U700 ( .A1(grant[1]), .A2(dbg_uart_wishbone_dat_w[24]), .B1(n395), 
        .B2(mgmtsoc_dbus_dbus_dat_w[24]), .ZN(n5083) );
  inv0d0 U701 ( .I(n5083), .ZN(mprj_dat_o[24]) );
  aoi22d1 U702 ( .A1(n396), .A2(dbg_uart_wishbone_dat_w[10]), .B1(n1888), .B2(
        mgmtsoc_dbus_dbus_dat_w[10]), .ZN(n5068) );
  inv0d0 U703 ( .I(n5068), .ZN(mprj_dat_o[10]) );
  aoi22d1 U704 ( .A1(n396), .A2(dbg_uart_wishbone_dat_w[8]), .B1(n1888), .B2(
        mgmtsoc_dbus_dbus_dat_w[8]), .ZN(n5066) );
  inv0d0 U705 ( .I(n5066), .ZN(mprj_dat_o[8]) );
  aoi22d1 U706 ( .A1(n397), .A2(dbg_uart_wishbone_dat_w[14]), .B1(n395), .B2(
        mgmtsoc_dbus_dbus_dat_w[14]), .ZN(n5072) );
  inv0d0 U707 ( .I(n5072), .ZN(mprj_dat_o[14]) );
  aoi22d1 U708 ( .A1(n397), .A2(dbg_uart_wishbone_dat_w[15]), .B1(n395), .B2(
        mgmtsoc_dbus_dbus_dat_w[15]), .ZN(n5073) );
  inv0d0 U709 ( .I(n5073), .ZN(mprj_dat_o[15]) );
  aoi22d1 U710 ( .A1(n396), .A2(dbg_uart_wishbone_dat_w[11]), .B1(n1888), .B2(
        mgmtsoc_dbus_dbus_dat_w[11]), .ZN(n5069) );
  inv0d0 U711 ( .I(n5069), .ZN(mprj_dat_o[11]) );
  aoi22d1 U712 ( .A1(n396), .A2(dbg_uart_wishbone_dat_w[31]), .B1(n395), .B2(
        mgmtsoc_dbus_dbus_dat_w[31]), .ZN(n5092) );
  inv0d0 U713 ( .I(n5092), .ZN(mprj_dat_o[31]) );
  aoi22d1 U714 ( .A1(n397), .A2(dbg_uart_wishbone_dat_w[21]), .B1(n1888), .B2(
        mgmtsoc_dbus_dbus_dat_w[21]), .ZN(n5080) );
  inv0d0 U715 ( .I(n5080), .ZN(mprj_dat_o[21]) );
  aoi22d1 U716 ( .A1(grant[1]), .A2(dbg_uart_wishbone_dat_w[25]), .B1(n395), 
        .B2(mgmtsoc_dbus_dbus_dat_w[25]), .ZN(n5084) );
  inv0d0 U717 ( .I(n5084), .ZN(mprj_dat_o[25]) );
  aoi22d1 U718 ( .A1(grant[1]), .A2(dbg_uart_wishbone_dat_w[30]), .B1(n395), 
        .B2(mgmtsoc_dbus_dbus_dat_w[30]), .ZN(n5091) );
  inv0d0 U719 ( .I(n5091), .ZN(mprj_dat_o[30]) );
  aoi22d1 U720 ( .A1(grant[1]), .A2(dbg_uart_wishbone_dat_w[23]), .B1(n395), 
        .B2(mgmtsoc_dbus_dbus_dat_w[23]), .ZN(n5082) );
  inv0d0 U721 ( .I(n5082), .ZN(mprj_dat_o[23]) );
  aoi22d1 U722 ( .A1(grant[1]), .A2(dbg_uart_wishbone_dat_w[27]), .B1(n394), 
        .B2(mgmtsoc_dbus_dbus_dat_w[27]), .ZN(n5087) );
  inv0d0 U723 ( .I(n5087), .ZN(mprj_dat_o[27]) );
  aoi22d1 U724 ( .A1(n397), .A2(dbg_uart_wishbone_dat_w[20]), .B1(n394), .B2(
        mgmtsoc_dbus_dbus_dat_w[20]), .ZN(n5079) );
  inv0d0 U725 ( .I(n5079), .ZN(mprj_dat_o[20]) );
  aoi22d1 U726 ( .A1(grant[1]), .A2(dbg_uart_wishbone_dat_w[28]), .B1(n394), 
        .B2(mgmtsoc_dbus_dbus_dat_w[28]), .ZN(n5088) );
  inv0d0 U727 ( .I(n5088), .ZN(mprj_dat_o[28]) );
  aoi22d1 U728 ( .A1(n397), .A2(dbg_uart_wishbone_dat_w[17]), .B1(n395), .B2(
        mgmtsoc_dbus_dbus_dat_w[17]), .ZN(n5075) );
  inv0d0 U729 ( .I(n5075), .ZN(mprj_dat_o[17]) );
  aoi22d1 U730 ( .A1(grant[1]), .A2(dbg_uart_wishbone_dat_w[29]), .B1(n394), 
        .B2(mgmtsoc_dbus_dbus_dat_w[29]), .ZN(n5090) );
  inv0d0 U731 ( .I(n5090), .ZN(mprj_dat_o[29]) );
  aoi22d1 U732 ( .A1(n397), .A2(dbg_uart_wishbone_dat_w[16]), .B1(n395), .B2(
        mgmtsoc_dbus_dbus_dat_w[16]), .ZN(n5074) );
  inv0d0 U733 ( .I(n5074), .ZN(mprj_dat_o[16]) );
  aoi22d1 U734 ( .A1(n397), .A2(dbg_uart_wishbone_dat_w[19]), .B1(n395), .B2(
        mgmtsoc_dbus_dbus_dat_w[19]), .ZN(n5078) );
  inv0d0 U735 ( .I(n5078), .ZN(mprj_dat_o[19]) );
  aoi22d1 U736 ( .A1(n397), .A2(dbg_uart_wishbone_dat_w[18]), .B1(n1888), .B2(
        mgmtsoc_dbus_dbus_dat_w[18]), .ZN(n5076) );
  inv0d0 U737 ( .I(n5076), .ZN(mprj_dat_o[18]) );
  aoi22d1 U738 ( .A1(n396), .A2(dbg_uart_wishbone_dat_w[12]), .B1(n395), .B2(
        mgmtsoc_dbus_dbus_dat_w[12]), .ZN(n5070) );
  inv0d0 U739 ( .I(n5070), .ZN(mprj_dat_o[12]) );
  aoi22d1 U740 ( .A1(n396), .A2(dbg_uart_wishbone_dat_w[9]), .B1(n395), .B2(
        mgmtsoc_dbus_dbus_dat_w[9]), .ZN(n5067) );
  inv0d0 U741 ( .I(n5067), .ZN(mprj_dat_o[9]) );
  aoi22d1 U742 ( .A1(n397), .A2(dbg_uart_wishbone_dat_w[13]), .B1(n395), .B2(
        mgmtsoc_dbus_dbus_dat_w[13]), .ZN(n5071) );
  inv0d0 U743 ( .I(n5071), .ZN(mprj_dat_o[13]) );
  aoi211d1 U744 ( .C1(csrbank0_reset0_w[0]), .C2(mgmtsoc_reset_re), .A(
        mgmtsoc_vexriscv_debug_reset), .B(csrbank0_reset0_w[1]), .ZN(n398) );
  nd02d1 U745 ( .A1(n398), .A2(n5301), .ZN(_2_net_) );
  buffd1 U746 ( .I(n6121), .Z(n6075) );
  buffd1 U747 ( .I(n6075), .Z(n6098) );
  buffd1 U748 ( .I(n6098), .Z(n6032) );
  buffd1 U749 ( .I(n6032), .Z(n6115) );
  buffd1 U750 ( .I(n6115), .Z(n6052) );
  buffd1 U751 ( .I(n6052), .Z(n6053) );
  buffd1 U752 ( .I(n6128), .Z(n6023) );
  buffd1 U753 ( .I(n6023), .Z(n6118) );
  buffd1 U754 ( .I(n6118), .Z(n6119) );
  buffd1 U755 ( .I(n6119), .Z(n6120) );
  buffd1 U756 ( .I(n6120), .Z(n6117) );
  buffd1 U757 ( .I(n6117), .Z(n6031) );
  buffd1 U758 ( .I(n6031), .Z(n6030) );
  buffd1 U759 ( .I(n6075), .Z(n6055) );
  buffd1 U760 ( .I(n6100), .Z(n6125) );
  buffd1 U761 ( .I(n6125), .Z(n6046) );
  buffd1 U762 ( .I(n6121), .Z(n6084) );
  buffd1 U763 ( .I(n6084), .Z(n6124) );
  buffd1 U764 ( .I(n6124), .Z(n6102) );
  buffd1 U765 ( .I(n6102), .Z(n6127) );
  buffd1 U766 ( .I(n6115), .Z(n6050) );
  buffd1 U767 ( .I(n6121), .Z(n6076) );
  buffd1 U768 ( .I(n6076), .Z(n6097) );
  buffd1 U769 ( .I(n6097), .Z(n6126) );
  buffd1 U770 ( .I(n6126), .Z(n6035) );
  buffd1 U771 ( .I(n6125), .Z(n6087) );
  buffd1 U772 ( .I(n6087), .Z(n6113) );
  buffd1 U773 ( .I(n6113), .Z(n6040) );
  buffd1 U774 ( .I(n6040), .Z(n6027) );
  buffd1 U775 ( .I(n6115), .Z(n6034) );
  buffd1 U776 ( .I(n6121), .Z(n6074) );
  buffd1 U777 ( .I(n6074), .Z(n6099) );
  buffd1 U778 ( .I(n6099), .Z(n6028) );
  buffd1 U779 ( .I(n6118), .Z(n6064) );
  buffd1 U780 ( .I(n6118), .Z(n6065) );
  buffd1 U781 ( .I(n6105), .Z(n6081) );
  buffd1 U782 ( .I(n6118), .Z(n6063) );
  buffd1 U783 ( .I(n6023), .Z(n6116) );
  buffd1 U784 ( .I(n6116), .Z(n6062) );
  buffd1 U785 ( .I(n6062), .Z(n6056) );
  buffd1 U786 ( .I(n6120), .Z(n6072) );
  buffd1 U787 ( .I(n6120), .Z(n6073) );
  buffd1 U788 ( .I(n6120), .Z(n6071) );
  buffd1 U789 ( .I(n6121), .Z(n6086) );
  buffd1 U790 ( .I(n6116), .Z(n6058) );
  buffd1 U791 ( .I(n6058), .Z(n6104) );
  buffd1 U792 ( .I(n6120), .Z(n6069) );
  buffd1 U793 ( .I(n6117), .Z(n6066) );
  buffd1 U794 ( .I(n6117), .Z(n6068) );
  buffd1 U795 ( .I(n6118), .Z(n6067) );
  buffd1 U796 ( .I(n6120), .Z(n6070) );
  buffd1 U797 ( .I(n6098), .Z(n6022) );
  buffd1 U798 ( .I(n6022), .Z(n6051) );
  buffd1 U799 ( .I(n6047), .Z(n6048) );
  buffd1 U800 ( .I(n6113), .Z(n6049) );
  buffd1 U801 ( .I(n6113), .Z(n6042) );
  buffd1 U802 ( .I(n6113), .Z(n6043) );
  buffd1 U803 ( .I(n6100), .Z(n6033) );
  buffd1 U804 ( .I(n6033), .Z(n6079) );
  buffd1 U805 ( .I(n6079), .Z(n6082) );
  buffd1 U806 ( .I(n6122), .Z(n6083) );
  buffd1 U807 ( .I(n6128), .Z(n6025) );
  buffd1 U808 ( .I(n6124), .Z(n6096) );
  buffd1 U809 ( .I(n6124), .Z(n6095) );
  buffd1 U810 ( .I(n6124), .Z(n6092) );
  buffd1 U811 ( .I(n6125), .Z(n6088) );
  buffd1 U812 ( .I(n6088), .Z(n6089) );
  buffd1 U813 ( .I(n6089), .Z(n6044) );
  buffd1 U814 ( .I(n6129), .Z(n6109) );
  buffd1 U815 ( .I(n6109), .Z(n6107) );
  buffd1 U816 ( .I(n6105), .Z(n6080) );
  buffd1 U817 ( .I(n6080), .Z(n6103) );
  buffd1 U818 ( .I(n6103), .Z(n6108) );
  buffd1 U819 ( .I(n6121), .Z(n6077) );
  buffd1 U820 ( .I(n6124), .Z(n6093) );
  buffd1 U821 ( .I(n6123), .Z(n6078) );
  buffd1 U822 ( .I(n6047), .Z(n6041) );
  buffd1 U823 ( .I(n6088), .Z(n6045) );
  buffd1 U824 ( .I(n6128), .Z(n6026) );
  buffd1 U825 ( .I(n6128), .Z(n6029) );
  buffd1 U826 ( .I(n6128), .Z(n6024) );
  buffd1 U827 ( .I(n6024), .Z(n6057) );
  buffd1 U828 ( .I(n6128), .Z(n6112) );
  buffd1 U829 ( .I(n6112), .Z(n6094) );
  buffd1 U830 ( .I(n6116), .Z(n6060) );
  buffd1 U831 ( .I(n6060), .Z(n6061) );
  buffd1 U832 ( .I(n6061), .Z(n6059) );
  buffd1 U833 ( .I(n6059), .Z(n6054) );
  buffd1 U834 ( .I(n6054), .Z(n6091) );
  buffd1 U835 ( .I(n6112), .Z(n6090) );
  buffd1 U836 ( .I(n6047), .Z(n6114) );
  buffd1 U837 ( .I(n6114), .Z(n6037) );
  buffd1 U838 ( .I(n6037), .Z(n6038) );
  buffd1 U839 ( .I(n6114), .Z(n6036) );
  buffd1 U840 ( .I(n6036), .Z(n6106) );
  buffd1 U841 ( .I(n6037), .Z(n6039) );
  inv0d0 U842 ( .I(uart_phy_tx_phase[11]), .ZN(n673) );
  inv0d0 U843 ( .I(uart_phy_tx_phase[9]), .ZN(n1463) );
  inv0d0 U844 ( .I(n1464), .ZN(n1465) );
  nd02d0 U845 ( .A1(n1463), .A2(n1465), .ZN(n1009) );
  inv0d0 U846 ( .I(n674), .ZN(n675) );
  nd02d0 U847 ( .A1(n673), .A2(n675), .ZN(n1028) );
  inv0d0 U848 ( .I(n1030), .ZN(n399) );
  aoim22d1 U849 ( .A1(uart_phy_tx_phase[13]), .A2(n399), .B1(n399), .B2(
        uart_phy_tx_phase[13]), .Z(n400) );
  inv0d0 U850 ( .I(rs232phy_rs232phytx_state), .ZN(n2848) );
  inv0d1 U851 ( .I(n2848), .ZN(n2868) );
  nd12d0 U852 ( .A1(n400), .A2(n2868), .ZN(N3585) );
  nr04d0 U853 ( .A1(dbg_uart_count[17]), .A2(dbg_uart_count[19]), .A3(
        dbg_uart_count[18]), .A4(dbg_uart_count[2]), .ZN(n404) );
  nr04d0 U854 ( .A1(dbg_uart_count[9]), .A2(dbg_uart_count[4]), .A3(
        dbg_uart_count[5]), .A4(dbg_uart_count[0]), .ZN(n403) );
  nr04d0 U855 ( .A1(dbg_uart_count[10]), .A2(dbg_uart_count[8]), .A3(
        dbg_uart_count[12]), .A4(dbg_uart_count[3]), .ZN(n402) );
  nr04d0 U856 ( .A1(dbg_uart_count[11]), .A2(dbg_uart_count[6]), .A3(
        dbg_uart_count[7]), .A4(dbg_uart_count[1]), .ZN(n401) );
  nr04d0 U857 ( .A1(dbg_uart_count[15]), .A2(dbg_uart_count[13]), .A3(
        dbg_uart_count[14]), .A4(dbg_uart_count[16]), .ZN(n405) );
  nd02d0 U858 ( .A1(n5955), .A2(n2497), .ZN(n2504) );
  nd02d0 U859 ( .A1(uartwishbonebridge_state[1]), .A2(
        uartwishbonebridge_state[2]), .ZN(n408) );
  inv0d0 U860 ( .I(uartwishbonebridge_state[2]), .ZN(n407) );
  nd02d0 U861 ( .A1(n5296), .A2(n407), .ZN(n1514) );
  aoi22d1 U862 ( .A1(uartwishbonebridge_state[0]), .A2(n408), .B1(n1514), .B2(
        n5488), .ZN(n2482) );
  nr02d1 U863 ( .A1(n2504), .A2(n2482), .ZN(n1171) );
  inv0d0 U864 ( .I(n1171), .ZN(n409) );
  nr02d0 U865 ( .A1(dbg_uart_count[0]), .A2(n409), .ZN(n4088) );
  inv0d0 U866 ( .I(litespiphy_state[0]), .ZN(n1544) );
  nr02d0 U867 ( .A1(litespiphy_state[1]), .A2(n1544), .ZN(n4857) );
  inv0d0 U868 ( .I(n4857), .ZN(n5732) );
  inv0d0 U869 ( .I(mgmtsoc_litespisdrphycore_div[5]), .ZN(n4868) );
  inv0d0 U870 ( .I(mgmtsoc_litespisdrphycore_div[6]), .ZN(n4869) );
  aoi22d1 U871 ( .A1(mgmtsoc_litespisdrphycore_cnt[5]), .A2(n4868), .B1(
        mgmtsoc_litespisdrphycore_cnt[6]), .B2(n4869), .ZN(n535) );
  inv0d0 U872 ( .I(mgmtsoc_litespisdrphycore_div[4]), .ZN(n4867) );
  inv0d0 U873 ( .I(mgmtsoc_litespisdrphycore_div[2]), .ZN(n4864) );
  inv0d0 U874 ( .I(mgmtsoc_litespisdrphycore_div[1]), .ZN(n4863) );
  aoi22d1 U875 ( .A1(mgmtsoc_litespisdrphycore_cnt[2]), .A2(n4864), .B1(
        mgmtsoc_litespisdrphycore_cnt[1]), .B2(n4863), .ZN(n526) );
  inv0d0 U876 ( .I(mgmtsoc_litespisdrphycore_div[0]), .ZN(n665) );
  oai22d1 U877 ( .A1(mgmtsoc_litespisdrphycore_cnt[1]), .A2(n4863), .B1(
        mgmtsoc_litespisdrphycore_cnt[0]), .B2(n665), .ZN(n530) );
  inv0d0 U878 ( .I(mgmtsoc_litespisdrphycore_div[3]), .ZN(n4865) );
  oai22d1 U879 ( .A1(mgmtsoc_litespisdrphycore_cnt[3]), .A2(n4865), .B1(
        mgmtsoc_litespisdrphycore_cnt[2]), .B2(n4864), .ZN(n528) );
  nd02d0 U880 ( .A1(mgmtsoc_litespisdrphycore_cnt[3]), .A2(n4865), .ZN(n410)
         );
  aon211d1 U881 ( .C1(n526), .C2(n530), .B(n528), .A(n410), .ZN(n412) );
  oai22d1 U882 ( .A1(mgmtsoc_litespisdrphycore_cnt[4]), .A2(n4867), .B1(
        mgmtsoc_litespisdrphycore_cnt[5]), .B2(n4868), .ZN(n529) );
  inv0d0 U883 ( .I(n529), .ZN(n411) );
  aon211d1 U884 ( .C1(mgmtsoc_litespisdrphycore_cnt[4]), .C2(n4867), .B(n412), 
        .A(n411), .ZN(n414) );
  inv0d0 U885 ( .I(mgmtsoc_litespisdrphycore_div[7]), .ZN(n4872) );
  oai22d1 U886 ( .A1(mgmtsoc_litespisdrphycore_cnt[6]), .A2(n4869), .B1(
        mgmtsoc_litespisdrphycore_cnt[7]), .B2(n4872), .ZN(n531) );
  nd02d0 U887 ( .A1(mgmtsoc_litespisdrphycore_cnt[7]), .A2(n4872), .ZN(n413)
         );
  aon211d1 U888 ( .C1(n535), .C2(n414), .B(n531), .A(n413), .ZN(n4859) );
  inv0d0 U889 ( .I(n993), .ZN(n415) );
  nr02d0 U890 ( .A1(mgmtsoc_litespisdrphycore_cnt[0]), .A2(n415), .ZN(N5443)
         );
  nr02d0 U891 ( .A1(spimaster_state[0]), .A2(spimaster_state[1]), .ZN(n3085)
         );
  nr04d0 U892 ( .A1(spi_master_clk_divider0[3]), .A2(
        spi_master_clk_divider0[2]), .A3(spi_master_clk_divider0[1]), .A4(
        spi_master_clk_divider0[0]), .ZN(n422) );
  inv0d0 U893 ( .I(spi_master_clk_divider0[4]), .ZN(n3067) );
  nd02d0 U894 ( .A1(n422), .A2(n3067), .ZN(n438) );
  nr02d0 U895 ( .A1(spi_master_clk_divider0[5]), .A2(n438), .ZN(n420) );
  inv0d0 U896 ( .I(spi_master_clk_divider0[6]), .ZN(n493) );
  nd02d0 U897 ( .A1(n420), .A2(n493), .ZN(n439) );
  nr02d0 U898 ( .A1(spi_master_clk_divider0[7]), .A2(n439), .ZN(n428) );
  inv0d0 U899 ( .I(spi_master_clk_divider0[8]), .ZN(n3072) );
  mx02d1 U900 ( .I0(n3072), .I1(spi_master_clk_divider0[8]), .S(
        spi_master_clk_divider1[8]), .Z(n427) );
  inv0d0 U901 ( .I(spi_master_clk_divider0[2]), .ZN(n3065) );
  mx02d1 U902 ( .I0(n3065), .I1(spi_master_clk_divider0[2]), .S(
        spi_master_clk_divider1[2]), .Z(n418) );
  nr02d0 U903 ( .A1(spi_master_clk_divider0[1]), .A2(
        spi_master_clk_divider0[0]), .ZN(n417) );
  oai22d1 U904 ( .A1(n417), .A2(n418), .B1(spi_master_clk_divider0[0]), .B2(
        spi_master_clk_divider1[0]), .ZN(n416) );
  aoi221d1 U905 ( .B1(n418), .B2(n417), .C1(spi_master_clk_divider0[0]), .C2(
        spi_master_clk_divider1[0]), .A(n416), .ZN(n425) );
  mx02d1 U906 ( .I0(n3067), .I1(spi_master_clk_divider0[4]), .S(
        spi_master_clk_divider1[4]), .Z(n423) );
  mx02d1 U907 ( .I0(n493), .I1(spi_master_clk_divider0[6]), .S(
        spi_master_clk_divider1[6]), .Z(n421) );
  oai22d1 U908 ( .A1(n422), .A2(n423), .B1(n421), .B2(n420), .ZN(n419) );
  aoi221d1 U909 ( .B1(n423), .B2(n422), .C1(n421), .C2(n420), .A(n419), .ZN(
        n424) );
  oai211d1 U910 ( .C1(n428), .C2(n427), .A(n425), .B(n424), .ZN(n426) );
  aoi21d1 U911 ( .B1(n428), .B2(n427), .A(n426), .ZN(n459) );
  inv0d0 U912 ( .I(spi_master_clk_divider0[10]), .ZN(n3074) );
  mx02d1 U913 ( .I0(n3074), .I1(spi_master_clk_divider0[10]), .S(
        spi_master_clk_divider1[10]), .Z(n432) );
  nd02d0 U914 ( .A1(n428), .A2(n3072), .ZN(n433) );
  nr02d0 U915 ( .A1(spi_master_clk_divider0[9]), .A2(n433), .ZN(n431) );
  inv0d0 U916 ( .I(spi_master_clk_divider0[12]), .ZN(n3076) );
  mx02d1 U917 ( .I0(n3076), .I1(spi_master_clk_divider0[12]), .S(
        spi_master_clk_divider1[12]), .Z(n430) );
  inv0d0 U918 ( .I(spi_master_clk_divider0[11]), .ZN(n3075) );
  an02d0 U919 ( .A1(n431), .A2(n3074), .Z(n454) );
  an02d0 U920 ( .A1(n3075), .A2(n454), .Z(n450) );
  oai22d1 U921 ( .A1(n450), .A2(n430), .B1(n431), .B2(n432), .ZN(n429) );
  aoi221d1 U922 ( .B1(n432), .B2(n431), .C1(n430), .C2(n450), .A(n429), .ZN(
        n458) );
  inv0d0 U923 ( .I(n433), .ZN(n449) );
  inv0d0 U924 ( .I(spi_master_clk_divider0[9]), .ZN(n3073) );
  mx02d1 U925 ( .I0(n3073), .I1(spi_master_clk_divider0[9]), .S(
        spi_master_clk_divider1[9]), .Z(n448) );
  inv0d0 U926 ( .I(spi_master_clk_divider0[3]), .ZN(n3066) );
  mx02d1 U927 ( .I0(n3066), .I1(spi_master_clk_divider0[3]), .S(
        spi_master_clk_divider1[3]), .Z(n437) );
  nr03d0 U928 ( .A1(spi_master_clk_divider0[2]), .A2(
        spi_master_clk_divider0[1]), .A3(spi_master_clk_divider0[0]), .ZN(n436) );
  aoim22d1 U929 ( .A1(spi_master_clk_divider0[1]), .A2(
        spi_master_clk_divider0[0]), .B1(spi_master_clk_divider0[0]), .B2(
        spi_master_clk_divider0[1]), .Z(n435) );
  oai22d1 U930 ( .A1(n436), .A2(n437), .B1(spi_master_clk_divider1[1]), .B2(
        n435), .ZN(n434) );
  aoi221d1 U931 ( .B1(n437), .B2(n436), .C1(spi_master_clk_divider1[1]), .C2(
        n435), .A(n434), .ZN(n446) );
  inv0d0 U932 ( .I(spi_master_clk_divider0[5]), .ZN(n3068) );
  mx02d1 U933 ( .I0(n3068), .I1(spi_master_clk_divider0[5]), .S(
        spi_master_clk_divider1[5]), .Z(n444) );
  inv0d0 U934 ( .I(n438), .ZN(n443) );
  inv0d0 U935 ( .I(spi_master_clk_divider0[7]), .ZN(n470) );
  mx02d1 U936 ( .I0(n470), .I1(spi_master_clk_divider0[7]), .S(
        spi_master_clk_divider1[7]), .Z(n442) );
  inv0d0 U937 ( .I(n439), .ZN(n441) );
  oai22d1 U938 ( .A1(n443), .A2(n444), .B1(n442), .B2(n441), .ZN(n440) );
  aoi221d1 U939 ( .B1(n444), .B2(n443), .C1(n442), .C2(n441), .A(n440), .ZN(
        n445) );
  oai211d1 U940 ( .C1(n449), .C2(n448), .A(n446), .B(n445), .ZN(n447) );
  aoi21d1 U941 ( .B1(n449), .B2(n448), .A(n447), .ZN(n457) );
  mx02d1 U942 ( .I0(n3075), .I1(spi_master_clk_divider0[11]), .S(
        spi_master_clk_divider1[11]), .Z(n455) );
  inv0d0 U943 ( .I(spi_master_clk_divider0[13]), .ZN(n3077) );
  mx02d1 U944 ( .I0(n3077), .I1(spi_master_clk_divider0[13]), .S(
        spi_master_clk_divider1[13]), .Z(n453) );
  nd02d0 U945 ( .A1(n3076), .A2(n450), .ZN(n460) );
  inv0d0 U946 ( .I(n460), .ZN(n452) );
  oai22d1 U947 ( .A1(n454), .A2(n455), .B1(n453), .B2(n452), .ZN(n451) );
  aoi221d1 U948 ( .B1(n455), .B2(n454), .C1(n453), .C2(n452), .A(n451), .ZN(
        n456) );
  nr02d0 U949 ( .A1(spi_master_clk_divider0[13]), .A2(n460), .ZN(n461) );
  inv0d0 U950 ( .I(spi_master_clk_divider0[14]), .ZN(n3078) );
  nd02d0 U951 ( .A1(n461), .A2(n3078), .ZN(n467) );
  nr02d0 U952 ( .A1(n461), .A2(n3078), .ZN(n462) );
  inv0d0 U953 ( .I(n462), .ZN(n466) );
  xr02d1 U954 ( .A1(spi_master_clk_divider0[15]), .A2(
        spi_master_clk_divider1[15]), .Z(n463) );
  nr02d0 U955 ( .A1(n462), .A2(n463), .ZN(n464) );
  aoi22d1 U956 ( .A1(spi_master_clk_divider1[14]), .A2(n464), .B1(n463), .B2(
        n467), .ZN(n465) );
  aon211d1 U957 ( .C1(n467), .C2(n466), .B(spi_master_clk_divider1[14]), .A(
        n465), .ZN(n468) );
  inv0d0 U958 ( .I(n1205), .ZN(n3089) );
  nr02d0 U959 ( .A1(spimaster_state[1]), .A2(n4677), .ZN(n1611) );
  nr04d0 U960 ( .A1(spi_master_clk_divider0[4]), .A2(
        spi_master_clk_divider0[3]), .A3(spi_master_clk_divider0[2]), .A4(
        spi_master_clk_divider0[1]), .ZN(n475) );
  nd02d0 U961 ( .A1(n475), .A2(n3068), .ZN(n494) );
  nr02d0 U962 ( .A1(spi_master_clk_divider0[6]), .A2(n494), .ZN(n472) );
  nd02d0 U963 ( .A1(n472), .A2(n470), .ZN(n495) );
  nr02d0 U964 ( .A1(spi_master_clk_divider0[8]), .A2(n495), .ZN(n483) );
  mx02d1 U965 ( .I0(n3073), .I1(spi_master_clk_divider0[9]), .S(
        spi_master_clk_divider1[8]), .Z(n482) );
  mx02d1 U966 ( .I0(n470), .I1(spi_master_clk_divider0[7]), .S(
        spi_master_clk_divider1[6]), .Z(n473) );
  oai22d1 U967 ( .A1(n472), .A2(n473), .B1(spi_master_clk_divider0[1]), .B2(
        spi_master_clk_divider1[0]), .ZN(n471) );
  aoi221d1 U968 ( .B1(n473), .B2(n472), .C1(spi_master_clk_divider0[1]), .C2(
        spi_master_clk_divider1[0]), .A(n471), .ZN(n480) );
  mx02d1 U969 ( .I0(n3066), .I1(spi_master_clk_divider0[3]), .S(
        spi_master_clk_divider1[2]), .Z(n478) );
  nr02d0 U970 ( .A1(spi_master_clk_divider0[2]), .A2(
        spi_master_clk_divider0[1]), .ZN(n477) );
  mx02d1 U971 ( .I0(n3068), .I1(spi_master_clk_divider0[5]), .S(
        spi_master_clk_divider1[4]), .Z(n476) );
  oai22d1 U972 ( .A1(n475), .A2(n476), .B1(n477), .B2(n478), .ZN(n474) );
  aoi221d1 U973 ( .B1(n478), .B2(n477), .C1(n476), .C2(n475), .A(n474), .ZN(
        n479) );
  oai211d1 U974 ( .C1(n483), .C2(n482), .A(n480), .B(n479), .ZN(n481) );
  aoi21d1 U975 ( .B1(n483), .B2(n482), .A(n481), .ZN(n515) );
  mx02d1 U976 ( .I0(n3075), .I1(spi_master_clk_divider0[11]), .S(
        spi_master_clk_divider1[10]), .Z(n487) );
  nd02d0 U977 ( .A1(n483), .A2(n3073), .ZN(n506) );
  nr02d0 U978 ( .A1(spi_master_clk_divider0[10]), .A2(n506), .ZN(n486) );
  mx02d1 U979 ( .I0(n3077), .I1(spi_master_clk_divider0[13]), .S(
        spi_master_clk_divider1[12]), .Z(n485) );
  an02d0 U980 ( .A1(n486), .A2(n3075), .Z(n508) );
  an02d0 U981 ( .A1(n3076), .A2(n508), .Z(n488) );
  oai22d1 U982 ( .A1(n486), .A2(n487), .B1(n485), .B2(n488), .ZN(n484) );
  aoi221d1 U983 ( .B1(n487), .B2(n486), .C1(n485), .C2(n488), .A(n484), .ZN(
        n514) );
  nd02d0 U984 ( .A1(n3077), .A2(n488), .ZN(n516) );
  inv0d0 U985 ( .I(n516), .ZN(n505) );
  mx02d1 U986 ( .I0(n3078), .I1(spi_master_clk_divider0[14]), .S(
        spi_master_clk_divider1[13]), .Z(n504) );
  mx02d1 U987 ( .I0(n3067), .I1(spi_master_clk_divider0[4]), .S(
        spi_master_clk_divider1[3]), .Z(n492) );
  nr03d0 U988 ( .A1(spi_master_clk_divider0[3]), .A2(
        spi_master_clk_divider0[2]), .A3(spi_master_clk_divider0[1]), .ZN(n491) );
  aoim22d1 U989 ( .A1(spi_master_clk_divider0[2]), .A2(
        spi_master_clk_divider0[1]), .B1(spi_master_clk_divider0[1]), .B2(
        spi_master_clk_divider0[2]), .Z(n490) );
  oai22d1 U990 ( .A1(n491), .A2(n492), .B1(spi_master_clk_divider1[1]), .B2(
        n490), .ZN(n489) );
  aoi221d1 U991 ( .B1(n492), .B2(n491), .C1(spi_master_clk_divider1[1]), .C2(
        n490), .A(n489), .ZN(n502) );
  mx02d1 U992 ( .I0(n493), .I1(spi_master_clk_divider0[6]), .S(
        spi_master_clk_divider1[5]), .Z(n500) );
  inv0d0 U993 ( .I(n494), .ZN(n499) );
  mx02d1 U994 ( .I0(n3072), .I1(spi_master_clk_divider0[8]), .S(
        spi_master_clk_divider1[7]), .Z(n498) );
  inv0d0 U995 ( .I(n495), .ZN(n497) );
  oai22d1 U996 ( .A1(n499), .A2(n500), .B1(n498), .B2(n497), .ZN(n496) );
  aoi221d1 U997 ( .B1(n500), .B2(n499), .C1(n498), .C2(n497), .A(n496), .ZN(
        n501) );
  oai211d1 U998 ( .C1(n505), .C2(n504), .A(n502), .B(n501), .ZN(n503) );
  aoi21d1 U999 ( .B1(n505), .B2(n504), .A(n503), .ZN(n513) );
  mx02d1 U1000 ( .I0(n3074), .I1(spi_master_clk_divider0[10]), .S(
        spi_master_clk_divider1[9]), .Z(n511) );
  inv0d0 U1001 ( .I(n506), .ZN(n510) );
  mx02d1 U1002 ( .I0(n3076), .I1(spi_master_clk_divider0[12]), .S(
        spi_master_clk_divider1[11]), .Z(n509) );
  oai22d1 U1003 ( .A1(n510), .A2(n511), .B1(n509), .B2(n508), .ZN(n507) );
  aoi221d1 U1004 ( .B1(n511), .B2(n510), .C1(n509), .C2(n508), .A(n507), .ZN(
        n512) );
  nr02d0 U1005 ( .A1(spi_master_clk_divider0[14]), .A2(n516), .ZN(n517) );
  inv0d0 U1006 ( .I(spi_master_clk_divider0[15]), .ZN(n3079) );
  nd02d0 U1007 ( .A1(n517), .A2(n3079), .ZN(n522) );
  nr02d0 U1008 ( .A1(n517), .A2(n3079), .ZN(n518) );
  inv0d0 U1009 ( .I(n518), .ZN(n521) );
  nr02d0 U1010 ( .A1(n518), .A2(spi_master_clk_divider1[15]), .ZN(n519) );
  aoi22d1 U1011 ( .A1(spi_master_clk_divider1[14]), .A2(n519), .B1(
        spi_master_clk_divider1[15]), .B2(n522), .ZN(n520) );
  aon211d1 U1012 ( .C1(n522), .C2(n521), .B(spi_master_clk_divider1[14]), .A(
        n520), .ZN(n523) );
  nr02d0 U1013 ( .A1(n524), .A2(n523), .ZN(n4679) );
  nd02d1 U1014 ( .A1(n5288), .A2(n4679), .ZN(n4682) );
  inv0d0 U1015 ( .I(spimaster_state[0]), .ZN(n4625) );
  inv0d0 U1016 ( .I(spimaster_state[1]), .ZN(n4627) );
  nr02d0 U1017 ( .A1(n4625), .A2(n4627), .ZN(n4622) );
  nd02d0 U1018 ( .A1(n5288), .A2(n4660), .ZN(n4661) );
  nr13d1 U1019 ( .A1(dff2_en), .A2(n4878), .A3(dff2_bus_ack), .ZN(N5433) );
  nr03d0 U1020 ( .A1(n5492), .A2(dff_bus_ack), .A3(n525), .ZN(N5432) );
  aoi22d1 U1021 ( .A1(mgmtsoc_litespisdrphycore_cnt[4]), .A2(n4867), .B1(
        mgmtsoc_litespisdrphycore_cnt[0]), .B2(n665), .ZN(n534) );
  oaim21d1 U1022 ( .B1(n4865), .B2(mgmtsoc_litespisdrphycore_cnt[3]), .A(n526), 
        .ZN(n527) );
  aoi211d1 U1023 ( .C1(mgmtsoc_litespisdrphycore_cnt[7]), .C2(n4872), .A(n5732), .B(n527), .ZN(n533) );
  nr04d0 U1024 ( .A1(n531), .A2(n530), .A3(n529), .A4(n528), .ZN(n532) );
  nd12d0 U1025 ( .A1(n1613), .A2(mgmtsoc_litespisdrphycore_clk), .ZN(n5926) );
  inv0d0 U1026 ( .I(mgmtsoc_port_master_user_port_sink_payload_width[1]), .ZN(
        n4766) );
  nr02d0 U1027 ( .A1(n4685), .A2(n4766), .ZN(n5913) );
  inv0d0 U1028 ( .I(mgmtsoc_port_master_user_port_sink_payload_width[0]), .ZN(
        n4765) );
  inv0d0 U1029 ( .I(mgmtsoc_port_master_user_port_sink_payload_width[2]), .ZN(
        n4768) );
  inv0d0 U1030 ( .I(n5932), .ZN(n5928) );
  nd02d0 U1031 ( .A1(litespi_tx_mux_sel), .A2(
        mgmtsoc_port_master_user_port_sink_payload_width[3]), .ZN(n1251) );
  nr02d1 U1032 ( .A1(n5926), .A2(n1867), .ZN(n5886) );
  buffd1 U1033 ( .I(n5886), .Z(n5897) );
  inv0d0 U1034 ( .I(n1251), .ZN(n5949) );
  inv0d0 U1035 ( .I(n5913), .ZN(n1249) );
  nr02d0 U1036 ( .A1(n5926), .A2(n1866), .ZN(n654) );
  buffd1 U1037 ( .I(n654), .Z(n5870) );
  aoi22d1 U1038 ( .A1(n5897), .A2(mgmtsoc_litespisdrphycore_sr_out[18]), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[12]), .ZN(n554) );
  inv0d0 U1039 ( .I(litespi_state[3]), .ZN(n1602) );
  nd02d0 U1040 ( .A1(litespi_state[0]), .A2(n1602), .ZN(n1551) );
  nr02d0 U1041 ( .A1(litespi_tx_mux_sel), .A2(n1551), .ZN(n1871) );
  aoi21d1 U1042 ( .B1(litespi_tx_mux_sel), .B2(
        mgmtsoc_port_master_user_port_sink_payload_width[0]), .A(n1871), .ZN(
        n5922) );
  or02d0 U1043 ( .A1(n5922), .A2(n5926), .Z(n5925) );
  nr04d0 U1044 ( .A1(n5932), .A2(n5913), .A3(n5949), .A4(n5925), .ZN(n5874) );
  inv0d0 U1045 ( .I(n5874), .ZN(n5908) );
  inv0d2 U1046 ( .I(n5908), .ZN(n5902) );
  inv0d0 U1047 ( .I(mgmtsoc_port_master_user_port_sink_payload_width[3]), .ZN(
        n4769) );
  nr02d1 U1048 ( .A1(n5926), .A2(n1870), .ZN(n5885) );
  buffd1 U1049 ( .I(n5885), .Z(n5893) );
  aoi22d1 U1050 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[19]), .B1(
        n5893), .B2(mgmtsoc_litespisdrphycore_sr_out[16]), .ZN(n553) );
  inv0d0 U1051 ( .I(n5926), .ZN(n1605) );
  nr04d0 U1052 ( .A1(mgmtsoc_litespisdrphycore_count[3]), .A2(
        mgmtsoc_litespisdrphycore_count[2]), .A3(
        mgmtsoc_litespisdrphycore_count[1]), .A4(
        mgmtsoc_litespisdrphycore_count[0]), .ZN(n4856) );
  aon211d1 U1053 ( .C1(litespi_tx_mux_sel), .C2(
        mgmtsoc_port_master_user_port_sink_valid), .B(n1871), .A(n4856), .ZN(
        n536) );
  nr03d1 U1054 ( .A1(litespiphy_state[0]), .A2(litespiphy_state[1]), .A3(n536), 
        .ZN(n5941) );
  aor211d1 U1055 ( .C1(n1605), .C2(n5735), .A(n5941), .B(n5874), .Z(n5906) );
  inv0d1 U1056 ( .I(n5906), .ZN(n5871) );
  inv0d0 U1057 ( .I(mgmtsoc_litespimmap_spi_dummy_bits[3]), .ZN(n4815) );
  inv0d0 U1058 ( .I(n1871), .ZN(n1595) );
  oan211d1 U1059 ( .C1(litespi_state[1]), .C2(n4815), .B(litespi_state[2]), 
        .A(n1595), .ZN(n537) );
  aoi21d1 U1060 ( .B1(litespi_tx_mux_sel), .B2(
        mgmtsoc_port_master_user_port_sink_payload_len[3]), .A(n537), .ZN(
        n5938) );
  inv0d0 U1061 ( .I(litespi_state[2]), .ZN(n543) );
  nr03d0 U1062 ( .A1(litespi_state[1]), .A2(n543), .A3(n1595), .ZN(n538) );
  inv0d0 U1063 ( .I(mgmtsoc_port_master_user_port_sink_payload_len[0]), .ZN(
        n4757) );
  nr02d1 U1064 ( .A1(n4685), .A2(n4757), .ZN(n5801) );
  buffd1 U1065 ( .I(n5801), .Z(n5787) );
  aoi21d1 U1066 ( .B1(mgmtsoc_litespimmap_spi_dummy_bits[0]), .B2(n538), .A(
        n5787), .ZN(n613) );
  aoi22d1 U1067 ( .A1(litespi_tx_mux_sel), .A2(
        mgmtsoc_port_master_user_port_sink_payload_len[1]), .B1(n538), .B2(
        mgmtsoc_litespimmap_spi_dummy_bits[1]), .ZN(n5912) );
  inv0d0 U1068 ( .I(n541), .ZN(n542) );
  aoi22d1 U1069 ( .A1(litespi_tx_mux_sel), .A2(
        mgmtsoc_port_master_user_port_sink_payload_len[2]), .B1(n538), .B2(
        mgmtsoc_litespimmap_spi_dummy_bits[2]), .ZN(n5931) );
  nd02d0 U1070 ( .A1(n542), .A2(n5931), .ZN(n540) );
  aoi21d1 U1071 ( .B1(n5938), .B2(n540), .A(n564), .ZN(n661) );
  aoi22d1 U1072 ( .A1(litespi_tx_mux_sel), .A2(
        mgmtsoc_port_master_user_port_sink_payload_len[4]), .B1(n538), .B2(
        mgmtsoc_litespimmap_spi_dummy_bits[4]), .ZN(n539) );
  nd03d0 U1073 ( .A1(n1871), .A2(litespi_state[1]), .A3(n543), .ZN(n1594) );
  nd02d0 U1074 ( .A1(n539), .A2(n1594), .ZN(n1252) );
  nr02d0 U1075 ( .A1(n1252), .A2(n5778), .ZN(n547) );
  aoi21d1 U1076 ( .B1(n1252), .B2(n5778), .A(n547), .ZN(n5785) );
  nr02d0 U1077 ( .A1(n659), .A2(n5785), .ZN(n685) );
  inv0d0 U1078 ( .I(n613), .ZN(n5921) );
  inv0d0 U1079 ( .I(n5912), .ZN(n612) );
  aoi21d1 U1080 ( .B1(n5921), .B2(n612), .A(n542), .ZN(n5821) );
  inv0d2 U1081 ( .I(n1594), .ZN(n621) );
  nr02d1 U1082 ( .A1(n4685), .A2(n5921), .ZN(n5800) );
  aoi222d1 U1083 ( .A1(mprj_adr_o[18]), .A2(n621), .B1(n5787), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[17]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[18]), .C2(n5800), .ZN(
        n604) );
  buffd1 U1084 ( .I(n5800), .Z(n5789) );
  aoi222d1 U1085 ( .A1(mprj_adr_o[20]), .A2(n621), .B1(n5801), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[19]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[20]), .C2(n5789), .ZN(
        n622) );
  inv0d1 U1086 ( .I(n5821), .ZN(n5818) );
  aoi22d1 U1087 ( .A1(n5821), .A2(n604), .B1(n622), .B2(n5818), .ZN(n5864) );
  inv0d1 U1088 ( .I(n5821), .ZN(n5804) );
  inv0d1 U1089 ( .I(n5804), .ZN(n5790) );
  aoi222d1 U1090 ( .A1(mprj_adr_o[14]), .A2(n621), .B1(n5787), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[13]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[14]), .C2(n5800), .ZN(
        n606) );
  aoi222d1 U1091 ( .A1(mprj_adr_o[16]), .A2(n621), .B1(n5787), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[15]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[16]), .C2(n5789), .ZN(
        n605) );
  aoi22d1 U1092 ( .A1(n5790), .A2(n606), .B1(n605), .B2(n5818), .ZN(n5861) );
  aoi22d1 U1093 ( .A1(n5862), .A2(n5864), .B1(n5861), .B2(n5830), .ZN(n688) );
  nd02d0 U1094 ( .A1(n1252), .A2(n659), .ZN(n689) );
  inv0d0 U1095 ( .I(n689), .ZN(n5783) );
  aoi222d1 U1096 ( .A1(mprj_adr_o[10]), .A2(n621), .B1(n5787), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[9]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[10]), .C2(n5789), .ZN(
        n608) );
  aoi222d1 U1097 ( .A1(mprj_adr_o[12]), .A2(n621), .B1(n5801), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[11]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[12]), .C2(n5789), .ZN(
        n607) );
  aoi22d1 U1098 ( .A1(n5821), .A2(n608), .B1(n607), .B2(n5818), .ZN(n5860) );
  aoi222d1 U1099 ( .A1(mprj_adr_o[6]), .A2(n621), .B1(n5787), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[5]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[6]), .C2(n5789), .ZN(
        n610) );
  aoi222d1 U1100 ( .A1(mprj_adr_o[8]), .A2(n621), .B1(n5787), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[7]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[8]), .C2(n5789), .ZN(
        n609) );
  aoi22d1 U1101 ( .A1(n5790), .A2(n610), .B1(n609), .B2(n5818), .ZN(n563) );
  aoi22d1 U1102 ( .A1(n5862), .A2(n5860), .B1(n563), .B2(n5830), .ZN(n578) );
  aoi22d1 U1103 ( .A1(n685), .A2(n688), .B1(n5783), .B2(n578), .ZN(n551) );
  nd02d0 U1104 ( .A1(n1871), .A2(n543), .ZN(n544) );
  inv0d0 U1105 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[0]), .ZN(
        n4725) );
  oai22d1 U1106 ( .A1(litespi_state[1]), .A2(n544), .B1(n4685), .B2(n4725), 
        .ZN(n5777) );
  inv0d0 U1107 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[2]), .ZN(
        n4727) );
  oai22d1 U1108 ( .A1(n5611), .A2(n1594), .B1(n4727), .B2(n4685), .ZN(n556) );
  inv0d0 U1109 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[1]), .ZN(
        n4726) );
  oai22d1 U1110 ( .A1(litespi_state[1]), .A2(n544), .B1(n4685), .B2(n4726), 
        .ZN(n555) );
  aoi22d1 U1111 ( .A1(n613), .A2(n556), .B1(n555), .B2(n5921), .ZN(n615) );
  aoi222d1 U1112 ( .A1(mprj_adr_o[4]), .A2(n621), .B1(n5801), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[3]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[4]), .C2(n5789), .ZN(
        n611) );
  aoi22d1 U1113 ( .A1(n5821), .A2(n615), .B1(n611), .B2(n5818), .ZN(n562) );
  aoi22d1 U1114 ( .A1(n545), .A2(n5777), .B1(n5862), .B2(n562), .ZN(n5896) );
  inv0d0 U1115 ( .I(mgmtsoc_port_master_user_port_sink_payload_len[5]), .ZN(
        n4764) );
  oai211d1 U1116 ( .C1(litespi_state[1]), .C2(
        mgmtsoc_litespimmap_spi_dummy_bits[5]), .A(n1871), .B(litespi_state[2]), .ZN(n546) );
  oai21d1 U1117 ( .B1(n4685), .B2(n4764), .A(n546), .ZN(n1262) );
  inv0d0 U1118 ( .I(n547), .ZN(n549) );
  oai21d1 U1119 ( .B1(n1262), .B2(n549), .A(n5941), .ZN(n548) );
  aoi21d1 U1120 ( .B1(n1262), .B2(n549), .A(n548), .ZN(n5784) );
  nd12d0 U1121 ( .A1(n5785), .A2(n5784), .ZN(n648) );
  oai21d1 U1122 ( .B1(n5896), .B2(n5786), .A(n648), .ZN(n550) );
  aoi22d1 U1123 ( .A1(n5871), .A2(mgmtsoc_litespisdrphycore_sr_out[20]), .B1(
        n551), .B2(n550), .ZN(n552) );
  aoi22d1 U1124 ( .A1(n5897), .A2(mgmtsoc_litespisdrphycore_sr_out[21]), .B1(
        n5893), .B2(mgmtsoc_litespisdrphycore_sr_out[19]), .ZN(n561) );
  aoi22d1 U1125 ( .A1(n5874), .A2(mgmtsoc_litespisdrphycore_sr_out[22]), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[15]), .ZN(n560) );
  aoi222d1 U1126 ( .A1(mprj_adr_o[21]), .A2(n621), .B1(n5801), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[20]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[21]), .C2(n5800), .ZN(
        n641) );
  aoi222d1 U1127 ( .A1(mprj_adr_o[23]), .A2(n621), .B1(n5801), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[22]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[23]), .C2(n5800), .ZN(
        n5820) );
  aoi22d1 U1128 ( .A1(n5790), .A2(n641), .B1(n5820), .B2(n5818), .ZN(n5831) );
  aoi222d1 U1129 ( .A1(mprj_adr_o[17]), .A2(n621), .B1(n5800), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[17]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[16]), .C2(n5787), .ZN(
        n590) );
  aoi222d1 U1130 ( .A1(mprj_adr_o[19]), .A2(n621), .B1(n5787), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[18]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[19]), .C2(n5800), .ZN(
        n642) );
  aoi22d1 U1131 ( .A1(n5790), .A2(n590), .B1(n642), .B2(n5804), .ZN(n569) );
  aoi22d1 U1132 ( .A1(n5862), .A2(n5831), .B1(n569), .B2(n5830), .ZN(n5793) );
  aoi222d1 U1133 ( .A1(mprj_adr_o[13]), .A2(n621), .B1(n5800), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[13]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[12]), .C2(n5787), .ZN(
        n592) );
  aoi222d1 U1134 ( .A1(mprj_adr_o[15]), .A2(n621), .B1(n5787), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[14]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[15]), .C2(n5800), .ZN(
        n591) );
  aoi22d1 U1135 ( .A1(n5821), .A2(n592), .B1(n591), .B2(n5804), .ZN(n568) );
  aoi222d1 U1136 ( .A1(mprj_adr_o[9]), .A2(n621), .B1(n5789), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[9]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[8]), .C2(n5801), .ZN(
        n594) );
  aoi222d1 U1137 ( .A1(mprj_adr_o[11]), .A2(n621), .B1(n5787), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[10]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[11]), .C2(n5789), .ZN(
        n593) );
  aoi22d1 U1138 ( .A1(n5790), .A2(n594), .B1(n593), .B2(n5818), .ZN(n571) );
  aoi22d1 U1139 ( .A1(n5862), .A2(n568), .B1(n571), .B2(n5830), .ZN(n586) );
  aoi22d1 U1140 ( .A1(n685), .A2(n5793), .B1(n5783), .B2(n586), .ZN(n558) );
  aoi222d1 U1141 ( .A1(mprj_adr_o[5]), .A2(n621), .B1(n5789), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[5]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[4]), .C2(n5787), .ZN(
        n596) );
  aoi222d1 U1142 ( .A1(mprj_adr_o[7]), .A2(n621), .B1(n5787), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[6]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[7]), .C2(n5789), .ZN(
        n595) );
  aoi22d1 U1143 ( .A1(n5790), .A2(n596), .B1(n595), .B2(n5818), .ZN(n570) );
  aoi22d1 U1144 ( .A1(n613), .A2(n555), .B1(n5777), .B2(n5921), .ZN(n598) );
  aoi222d1 U1145 ( .A1(n556), .A2(n5921), .B1(
        mgmtsoc_port_master_user_port_sink_payload_data[3]), .B2(n5789), .C1(
        mprj_adr_o[3]), .C2(n621), .ZN(n597) );
  aoi22d1 U1146 ( .A1(n5790), .A2(n598), .B1(n597), .B2(n5818), .ZN(n572) );
  aoi22d1 U1147 ( .A1(n5862), .A2(n570), .B1(n572), .B2(n5830), .ZN(n5884) );
  oai21d1 U1148 ( .B1(n5786), .B2(n5884), .A(n648), .ZN(n557) );
  aoi22d1 U1149 ( .A1(n5871), .A2(mgmtsoc_litespisdrphycore_sr_out[23]), .B1(
        n558), .B2(n557), .ZN(n559) );
  aoi22d1 U1150 ( .A1(n5886), .A2(mgmtsoc_litespisdrphycore_sr_out[6]), .B1(
        n654), .B2(mgmtsoc_litespisdrphycore_sr_out[0]), .ZN(n567) );
  aoi22d1 U1151 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[7]), .B1(
        n5893), .B2(mgmtsoc_litespisdrphycore_sr_out[4]), .ZN(n566) );
  inv0d0 U1152 ( .I(n648), .ZN(n5780) );
  inv0d0 U1153 ( .I(n5862), .ZN(n5863) );
  aoi22d1 U1154 ( .A1(n5862), .A2(n563), .B1(n562), .B2(n5863), .ZN(n5876) );
  oaim22d1 U1155 ( .A1(n659), .A2(n5876), .B1(n5777), .B2(n564), .ZN(n5869) );
  aoi22d1 U1156 ( .A1(n5871), .A2(mgmtsoc_litespisdrphycore_sr_out[8]), .B1(
        n5780), .B2(n5869), .ZN(n565) );
  aoi22d1 U1157 ( .A1(n5897), .A2(mgmtsoc_litespisdrphycore_sr_out[17]), .B1(
        n5885), .B2(mgmtsoc_litespisdrphycore_sr_out[15]), .ZN(n577) );
  aoi22d1 U1158 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[18]), .B1(
        n654), .B2(mgmtsoc_litespisdrphycore_sr_out[11]), .ZN(n576) );
  aoi22d1 U1159 ( .A1(n5862), .A2(n569), .B1(n568), .B2(n5830), .ZN(n5834) );
  aoi22d1 U1160 ( .A1(n5862), .A2(n571), .B1(n570), .B2(n5830), .ZN(n582) );
  aoi22d1 U1161 ( .A1(n685), .A2(n5834), .B1(n5783), .B2(n582), .ZN(n574) );
  oai21d1 U1162 ( .B1(n5900), .B2(n5786), .A(n648), .ZN(n573) );
  aoi22d1 U1163 ( .A1(n5871), .A2(mgmtsoc_litespisdrphycore_sr_out[19]), .B1(
        n574), .B2(n573), .ZN(n575) );
  aoi22d1 U1164 ( .A1(n5885), .A2(mgmtsoc_litespisdrphycore_sr_out[8]), .B1(
        n654), .B2(mgmtsoc_litespisdrphycore_sr_out[4]), .ZN(n581) );
  aoi22d1 U1165 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[11]), .B1(
        n5886), .B2(mgmtsoc_litespisdrphycore_sr_out[10]), .ZN(n580) );
  inv0d1 U1166 ( .I(n5906), .ZN(n5901) );
  aoi22d1 U1167 ( .A1(n661), .A2(n578), .B1(n5896), .B2(n659), .ZN(n693) );
  aoi22d1 U1168 ( .A1(n5901), .A2(mgmtsoc_litespisdrphycore_sr_out[12]), .B1(
        n693), .B2(n5780), .ZN(n579) );
  aoi22d1 U1169 ( .A1(n5886), .A2(mgmtsoc_litespisdrphycore_sr_out[9]), .B1(
        n654), .B2(mgmtsoc_litespisdrphycore_sr_out[3]), .ZN(n585) );
  aoi22d1 U1170 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[10]), .B1(
        n5893), .B2(mgmtsoc_litespisdrphycore_sr_out[7]), .ZN(n584) );
  aoi22d1 U1171 ( .A1(n661), .A2(n582), .B1(n5900), .B2(n659), .ZN(n5837) );
  aoi22d1 U1172 ( .A1(n5901), .A2(mgmtsoc_litespisdrphycore_sr_out[11]), .B1(
        n5780), .B2(n5837), .ZN(n583) );
  aoi22d1 U1173 ( .A1(n5897), .A2(mgmtsoc_litespisdrphycore_sr_out[13]), .B1(
        n5893), .B2(mgmtsoc_litespisdrphycore_sr_out[11]), .ZN(n589) );
  aoi22d1 U1174 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[14]), .B1(
        n654), .B2(mgmtsoc_litespisdrphycore_sr_out[7]), .ZN(n588) );
  aoi22d1 U1175 ( .A1(n661), .A2(n586), .B1(n5884), .B2(n659), .ZN(n5796) );
  aoi22d1 U1176 ( .A1(n5871), .A2(mgmtsoc_litespisdrphycore_sr_out[15]), .B1(
        n5780), .B2(n5796), .ZN(n587) );
  aoi22d1 U1177 ( .A1(n5897), .A2(mgmtsoc_litespisdrphycore_sr_out[15]), .B1(
        n5885), .B2(mgmtsoc_litespisdrphycore_sr_out[13]), .ZN(n603) );
  aoi22d1 U1178 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[16]), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[9]), .ZN(n602) );
  aoi22d1 U1179 ( .A1(n5821), .A2(n591), .B1(n590), .B2(n5818), .ZN(n643) );
  aoi22d1 U1180 ( .A1(n5821), .A2(n593), .B1(n592), .B2(n5804), .ZN(n645) );
  aoi22d1 U1181 ( .A1(n5862), .A2(n643), .B1(n645), .B2(n5863), .ZN(n5853) );
  aoi22d1 U1182 ( .A1(n5790), .A2(n595), .B1(n594), .B2(n5804), .ZN(n644) );
  aoi22d1 U1183 ( .A1(n5790), .A2(n597), .B1(n596), .B2(n5804), .ZN(n647) );
  aoi22d1 U1184 ( .A1(n5862), .A2(n644), .B1(n647), .B2(n5863), .ZN(n655) );
  aoi22d1 U1185 ( .A1(n685), .A2(n5853), .B1(n5783), .B2(n655), .ZN(n600) );
  nr02d0 U1186 ( .A1(n5790), .A2(n598), .ZN(n646) );
  oai21d1 U1187 ( .B1(n5911), .B2(n5786), .A(n648), .ZN(n599) );
  aoi22d1 U1188 ( .A1(n5871), .A2(mgmtsoc_litespisdrphycore_sr_out[17]), .B1(
        n600), .B2(n599), .ZN(n601) );
  aoi22d1 U1189 ( .A1(n5897), .A2(mgmtsoc_litespisdrphycore_sr_out[16]), .B1(
        n654), .B2(mgmtsoc_litespisdrphycore_sr_out[10]), .ZN(n620) );
  aoi22d1 U1190 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[17]), .B1(
        n5885), .B2(mgmtsoc_litespisdrphycore_sr_out[14]), .ZN(n619) );
  aoi22d1 U1191 ( .A1(n5821), .A2(n605), .B1(n604), .B2(n5804), .ZN(n623) );
  aoi22d1 U1192 ( .A1(n5790), .A2(n607), .B1(n606), .B2(n5804), .ZN(n625) );
  aoi22d1 U1193 ( .A1(n5862), .A2(n623), .B1(n625), .B2(n5863), .ZN(n5844) );
  aoi22d1 U1194 ( .A1(n5790), .A2(n609), .B1(n608), .B2(n5804), .ZN(n624) );
  aoi22d1 U1195 ( .A1(n5790), .A2(n611), .B1(n610), .B2(n5804), .ZN(n627) );
  aoi22d1 U1196 ( .A1(n5862), .A2(n624), .B1(n627), .B2(n5863), .ZN(n637) );
  aoi22d1 U1197 ( .A1(n685), .A2(n5844), .B1(n5783), .B2(n637), .ZN(n617) );
  oai21d1 U1198 ( .B1(n5790), .B2(n615), .A(n614), .ZN(n626) );
  oai21d1 U1199 ( .B1(n5905), .B2(n5786), .A(n648), .ZN(n616) );
  aoi22d1 U1200 ( .A1(n5871), .A2(mgmtsoc_litespisdrphycore_sr_out[18]), .B1(
        n617), .B2(n616), .ZN(n618) );
  aoi22d1 U1201 ( .A1(n5897), .A2(mgmtsoc_litespisdrphycore_sr_out[20]), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[14]), .ZN(n632) );
  aoi22d1 U1202 ( .A1(n5874), .A2(mgmtsoc_litespisdrphycore_sr_out[21]), .B1(
        n5893), .B2(mgmtsoc_litespisdrphycore_sr_out[18]), .ZN(n631) );
  aoi222d1 U1203 ( .A1(mprj_adr_o[22]), .A2(n621), .B1(n5801), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[21]), .C1(
        mgmtsoc_port_master_user_port_sink_payload_data[22]), .C2(n5789), .ZN(
        n686) );
  aoi22d1 U1204 ( .A1(n5790), .A2(n622), .B1(n686), .B2(n5804), .ZN(n5841) );
  aoi22d1 U1205 ( .A1(n5862), .A2(n5841), .B1(n623), .B2(n5830), .ZN(n5809) );
  aoi22d1 U1206 ( .A1(n5862), .A2(n625), .B1(n624), .B2(n5830), .ZN(n633) );
  aoi22d1 U1207 ( .A1(n685), .A2(n5809), .B1(n5783), .B2(n633), .ZN(n629) );
  aoi22d1 U1208 ( .A1(n5862), .A2(n627), .B1(n626), .B2(n5830), .ZN(n5889) );
  oai21d1 U1209 ( .B1(n5889), .B2(n5786), .A(n648), .ZN(n628) );
  aoi22d1 U1210 ( .A1(n5871), .A2(mgmtsoc_litespisdrphycore_sr_out[22]), .B1(
        n629), .B2(n628), .ZN(n630) );
  aoi22d1 U1211 ( .A1(n5897), .A2(mgmtsoc_litespisdrphycore_sr_out[12]), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[6]), .ZN(n636) );
  aoi22d1 U1212 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[13]), .B1(
        n5885), .B2(mgmtsoc_litespisdrphycore_sr_out[10]), .ZN(n635) );
  aoi22d1 U1213 ( .A1(n661), .A2(n633), .B1(n5889), .B2(n659), .ZN(n5812) );
  aoi22d1 U1214 ( .A1(n5871), .A2(mgmtsoc_litespisdrphycore_sr_out[14]), .B1(
        n5780), .B2(n5812), .ZN(n634) );
  aoi22d1 U1215 ( .A1(n5885), .A2(mgmtsoc_litespisdrphycore_sr_out[6]), .B1(
        n654), .B2(mgmtsoc_litespisdrphycore_sr_out[2]), .ZN(n640) );
  aoi22d1 U1216 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[9]), .B1(
        n5886), .B2(mgmtsoc_litespisdrphycore_sr_out[8]), .ZN(n639) );
  aoi22d1 U1217 ( .A1(n661), .A2(n637), .B1(n5905), .B2(n659), .ZN(n5847) );
  aoi22d1 U1218 ( .A1(n5871), .A2(mgmtsoc_litespisdrphycore_sr_out[10]), .B1(
        n5780), .B2(n5847), .ZN(n638) );
  aoi22d1 U1219 ( .A1(n5897), .A2(mgmtsoc_litespisdrphycore_sr_out[19]), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[13]), .ZN(n653) );
  aoi22d1 U1220 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[20]), .B1(
        n5893), .B2(mgmtsoc_litespisdrphycore_sr_out[17]), .ZN(n652) );
  aoi22d1 U1221 ( .A1(n5821), .A2(n642), .B1(n641), .B2(n5818), .ZN(n5850) );
  aoi22d1 U1222 ( .A1(n5862), .A2(n5850), .B1(n643), .B2(n5830), .ZN(n5824) );
  aoi22d1 U1223 ( .A1(n5862), .A2(n645), .B1(n644), .B2(n5830), .ZN(n660) );
  aoi22d1 U1224 ( .A1(n685), .A2(n5824), .B1(n5783), .B2(n660), .ZN(n650) );
  aoi22d1 U1225 ( .A1(n5862), .A2(n647), .B1(n646), .B2(n5830), .ZN(n5892) );
  oai21d1 U1226 ( .B1(n5892), .B2(n5786), .A(n648), .ZN(n649) );
  aoi22d1 U1227 ( .A1(n5871), .A2(mgmtsoc_litespisdrphycore_sr_out[21]), .B1(
        n650), .B2(n649), .ZN(n651) );
  aoi22d1 U1228 ( .A1(n5897), .A2(mgmtsoc_litespisdrphycore_sr_out[7]), .B1(
        n654), .B2(mgmtsoc_litespisdrphycore_sr_out[1]), .ZN(n658) );
  aoi22d1 U1229 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[8]), .B1(
        n5893), .B2(mgmtsoc_litespisdrphycore_sr_out[5]), .ZN(n657) );
  aoi22d1 U1230 ( .A1(n661), .A2(n655), .B1(n5911), .B2(n659), .ZN(n5856) );
  aoi22d1 U1231 ( .A1(n5901), .A2(mgmtsoc_litespisdrphycore_sr_out[9]), .B1(
        n5780), .B2(n5856), .ZN(n656) );
  aoi22d1 U1232 ( .A1(n5897), .A2(mgmtsoc_litespisdrphycore_sr_out[11]), .B1(
        n5885), .B2(mgmtsoc_litespisdrphycore_sr_out[9]), .ZN(n664) );
  aoi22d1 U1233 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[12]), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[5]), .ZN(n663) );
  aoi22d1 U1234 ( .A1(n661), .A2(n660), .B1(n5892), .B2(n659), .ZN(n5827) );
  aoi22d1 U1235 ( .A1(n5901), .A2(mgmtsoc_litespisdrphycore_sr_out[13]), .B1(
        n5780), .B2(n5827), .ZN(n662) );
  nr02d0 U1236 ( .A1(n665), .A2(n4860), .ZN(N4292) );
  nr02d0 U1237 ( .A1(n4869), .A2(n4860), .ZN(N4298) );
  nr02d0 U1238 ( .A1(n4863), .A2(n4860), .ZN(N4293) );
  nr02d0 U1239 ( .A1(n4872), .A2(n4860), .ZN(N4299) );
  nr02d0 U1240 ( .A1(n4868), .A2(n4860), .ZN(N4297) );
  inv0d0 U1241 ( .I(serial_rx), .ZN(n666) );
  nr02d0 U1242 ( .A1(debug_in), .A2(n666), .ZN(sys_uart_rx) );
  inv0d0 U1243 ( .I(csrbank16_mode0_w), .ZN(n667) );
  aoi22d1 U1244 ( .A1(csrbank16_mode0_w), .A2(gpioin3_gpioin3_in_pads_n_d), 
        .B1(csrbank16_edge0_w), .B2(n667), .ZN(n668) );
  mx02d1 U1245 ( .I0(csrbank16_in_w), .I1(n669), .S(n668), .Z(n1949) );
  nr02d0 U1246 ( .A1(n2516), .A2(n670), .ZN(N6236) );
  inv0d0 U1247 ( .I(csrbank18_in_w), .ZN(n672) );
  nr02d0 U1248 ( .A1(n2516), .A2(n1941), .ZN(N6239) );
  inv0d0 U1249 ( .I(csrbank18_mode0_w), .ZN(n1768) );
  aoi22d1 U1250 ( .A1(csrbank18_mode0_w), .A2(gpioin5_gpioin5_in_pads_n_d), 
        .B1(csrbank18_edge0_w), .B2(n1768), .ZN(n671) );
  mx02d1 U1251 ( .I0(csrbank18_in_w), .I1(n672), .S(n671), .Z(n1934) );
  aoi22d1 U1252 ( .A1(uart_phy_tx_phase[11]), .A2(n675), .B1(n674), .B2(n673), 
        .ZN(n676) );
  nd12d0 U1253 ( .A1(n676), .A2(n2868), .ZN(N3583) );
  inv0d0 U1254 ( .I(uart_phy_tx_phase[14]), .ZN(n678) );
  nr02d0 U1255 ( .A1(uart_phy_tx_phase[13]), .A2(n1030), .ZN(n677) );
  mx02d1 U1256 ( .I0(uart_phy_tx_phase[14]), .I1(n678), .S(n677), .Z(n679) );
  nd12d0 U1257 ( .A1(n679), .A2(n2868), .ZN(N3586) );
  inv0d0 U1258 ( .I(n680), .ZN(n681) );
  nr02d0 U1259 ( .A1(n2516), .A2(n1545), .ZN(N6301) );
  nr02d0 U1260 ( .A1(n2516), .A2(n683), .ZN(N6303) );
  inv0d0 U1261 ( .I(uart_phy_rx_phase[11]), .ZN(n1011) );
  inv0d0 U1262 ( .I(uart_phy_rx_phase[9]), .ZN(n1005) );
  inv0d0 U1263 ( .I(n1006), .ZN(n1007) );
  nd02d0 U1264 ( .A1(n1005), .A2(n1007), .ZN(n1015) );
  inv0d0 U1265 ( .I(n1012), .ZN(n1013) );
  nd02d0 U1266 ( .A1(n1011), .A2(n1013), .ZN(n1017) );
  nr03d0 U1267 ( .A1(uart_phy_rx_phase[14]), .A2(uart_phy_rx_phase[13]), .A3(
        n1022), .ZN(n1025) );
  inv0d0 U1268 ( .I(uart_phy_rx_phase[15]), .ZN(n1026) );
  nd02d0 U1269 ( .A1(n1025), .A2(n1026), .ZN(n1032) );
  nr03d0 U1270 ( .A1(uart_phy_rx_phase[18]), .A2(uart_phy_rx_phase[17]), .A3(
        n1037), .ZN(n1075) );
  nd12d0 U1271 ( .A1(uart_phy_rx_phase[19]), .A2(n1075), .ZN(n1108) );
  nr02d0 U1272 ( .A1(uart_phy_rx_phase[20]), .A2(n1108), .ZN(n1105) );
  inv0d0 U1273 ( .I(uart_phy_rx_phase[21]), .ZN(n1106) );
  nd02d0 U1274 ( .A1(n1105), .A2(n1106), .ZN(n1126) );
  nd12d0 U1275 ( .A1(n684), .A2(n1200), .ZN(N3670) );
  aoi22d1 U1276 ( .A1(n5886), .A2(mgmtsoc_litespisdrphycore_sr_out[26]), .B1(
        n5893), .B2(mgmtsoc_litespisdrphycore_sr_out[24]), .ZN(n697) );
  aoi22d1 U1277 ( .A1(n5874), .A2(mgmtsoc_litespisdrphycore_sr_out[27]), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[20]), .ZN(n696) );
  nd02d0 U1278 ( .A1(n5901), .A2(mgmtsoc_litespisdrphycore_sr_out[28]), .ZN(
        n695) );
  inv0d0 U1279 ( .I(n685), .ZN(n691) );
  aoi22d1 U1280 ( .A1(n5787), .A2(
        mgmtsoc_port_master_user_port_sink_payload_data[25]), .B1(n5789), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[26]), .ZN(n5805) );
  aoi22d1 U1281 ( .A1(n5801), .A2(
        mgmtsoc_port_master_user_port_sink_payload_data[27]), .B1(n5800), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[28]), .ZN(n5803) );
  aoi22d1 U1282 ( .A1(n5821), .A2(n5805), .B1(n5803), .B2(n5818), .ZN(n687) );
  aoi22d1 U1283 ( .A1(n5801), .A2(
        mgmtsoc_port_master_user_port_sink_payload_data[23]), .B1(n5789), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[24]), .ZN(n5806) );
  aoi22d1 U1284 ( .A1(n5821), .A2(n686), .B1(n5806), .B2(n5818), .ZN(n5865) );
  aoi22d1 U1285 ( .A1(n5862), .A2(n687), .B1(n5865), .B2(n5830), .ZN(n690) );
  oai22d1 U1286 ( .A1(n691), .A2(n690), .B1(n689), .B2(n688), .ZN(n692) );
  aon211d1 U1287 ( .C1(n5785), .C2(n693), .B(n692), .A(n5784), .ZN(n694) );
  nr03d0 U1288 ( .A1(count[2]), .A2(count[1]), .A3(count[0]), .ZN(n1288) );
  inv0d0 U1289 ( .I(n1288), .ZN(n698) );
  nr02d0 U1290 ( .A1(n698), .A2(count[3]), .ZN(n1286) );
  nr02d0 U1291 ( .A1(n1296), .A2(count[5]), .ZN(n701) );
  nr02d0 U1292 ( .A1(n1309), .A2(count[7]), .ZN(n1306) );
  nd12d0 U1293 ( .A1(count[8]), .A2(n1306), .ZN(n703) );
  inv0d0 U1294 ( .I(n703), .ZN(n699) );
  aoim22d1 U1295 ( .A1(count[9]), .A2(n699), .B1(n699), .B2(count[9]), .Z(n700) );
  nd12d0 U1296 ( .A1(n700), .A2(n1314), .ZN(n4526) );
  aoim22d1 U1297 ( .A1(count[6]), .A2(n701), .B1(n701), .B2(count[6]), .Z(n702) );
  nd12d0 U1298 ( .A1(n702), .A2(n1314), .ZN(n4523) );
  nr02d0 U1299 ( .A1(n703), .A2(count[9]), .ZN(n1311) );
  nd12d0 U1300 ( .A1(count[10]), .A2(n1311), .ZN(n1293) );
  nr02d0 U1301 ( .A1(n1293), .A2(count[11]), .ZN(n1290) );
  nd12d0 U1302 ( .A1(count[12]), .A2(n1290), .ZN(n1304) );
  nr02d0 U1303 ( .A1(n1304), .A2(count[13]), .ZN(n1283) );
  aoim22d1 U1304 ( .A1(count[14]), .A2(n1283), .B1(n1283), .B2(count[14]), .Z(
        n704) );
  nd12d0 U1305 ( .A1(n704), .A2(n1314), .ZN(n4531) );
  inv0d0 U1306 ( .I(n4579), .ZN(n1828) );
  inv0d0 U1307 ( .I(csrbank9_cs0_w[16]), .ZN(n4603) );
  nr02d0 U1308 ( .A1(n1828), .A2(n4603), .ZN(N4601) );
  inv0d0 U1309 ( .I(n6131), .ZN(n1979) );
  inv0d0 U1310 ( .I(n6132), .ZN(n1978) );
  inv0d0 U1311 ( .I(n6133), .ZN(n1977) );
  nr02d0 U1312 ( .A1(n1976), .A2(n1977), .ZN(N4995) );
  inv0d0 U1313 ( .I(n2654), .ZN(n2258) );
  nd02d0 U1314 ( .A1(n1944), .A2(n2258), .ZN(n1911) );
  nr02d0 U1315 ( .A1(n2516), .A2(n1911), .ZN(N6285) );
  inv0d0 U1316 ( .I(n1546), .ZN(n1597) );
  nd03d1 U1317 ( .A1(n1597), .A2(slave_sel_r[3]), .A3(n4685), .ZN(n5432) );
  inv0d2 U1318 ( .I(n5432), .ZN(n1459) );
  inv0d1 U1319 ( .I(n5425), .ZN(n5335) );
  aoi21d1 U1320 ( .B1(mgmtsoc_litespisdrphycore_source_payload_data[25]), .B2(
        n1459), .A(n5335), .ZN(n713) );
  buffd1 U1321 ( .I(slave_sel_r[0]), .Z(n5395) );
  aoi22d1 U1322 ( .A1(n5395), .A2(mgmtsoc_vexriscv_debug_bus_dat_r[1]), .B1(
        slave_sel_r[5]), .B2(hk_dat_i[1]), .ZN(n712) );
  nr04d0 U1323 ( .A1(interface9_bank_bus_dat_r[1]), .A2(
        interface10_bank_bus_dat_r[1]), .A3(interface11_bank_bus_dat_r[1]), 
        .A4(interface19_bank_bus_dat_r[1]), .ZN(n707) );
  nd02d1 U1324 ( .A1(state), .A2(slave_sel_r[6]), .ZN(n5356) );
  buffd1 U1325 ( .I(n5356), .Z(n5426) );
  buffd1 U1326 ( .I(slave_sel_r[4]), .Z(n5394) );
  buffd1 U1327 ( .I(slave_sel_r[2]), .Z(n5406) );
  aoi22d1 U1328 ( .A1(n5394), .A2(mprj_dat_i[1]), .B1(n5406), .B2(
        dff2_bus_dat_r[1]), .ZN(n705) );
  aon211d1 U1329 ( .C1(n707), .C2(n706), .B(n5426), .A(n705), .ZN(n708) );
  inv0d0 U1330 ( .I(n708), .ZN(n711) );
  inv0d0 U1331 ( .I(slave_sel_r[1]), .ZN(n709) );
  buffd1 U1332 ( .I(n5380), .Z(n5401) );
  nr02d1 U1333 ( .A1(mprj_adr_o[9]), .A2(n709), .ZN(n1409) );
  buffd1 U1334 ( .I(n1409), .Z(n5435) );
  aoi22d1 U1335 ( .A1(n5401), .A2(\RAM256/Do0_pre[1][1] ), .B1(n5435), .B2(
        \RAM256/Do0_pre[0][1] ), .ZN(n710) );
  aoi21d1 U1336 ( .B1(mgmtsoc_litespisdrphycore_source_payload_data[26]), .B2(
        n1459), .A(n5335), .ZN(n721) );
  buffd1 U1337 ( .I(slave_sel_r[5]), .Z(n5429) );
  aoi22d1 U1338 ( .A1(n5429), .A2(hk_dat_i[2]), .B1(n5406), .B2(
        dff2_bus_dat_r[2]), .ZN(n720) );
  nr04d0 U1339 ( .A1(interface9_bank_bus_dat_r[2]), .A2(
        interface10_bank_bus_dat_r[2]), .A3(interface11_bank_bus_dat_r[2]), 
        .A4(interface19_bank_bus_dat_r[2]), .ZN(n716) );
  nr04d0 U1340 ( .A1(interface0_bank_bus_dat_r[2]), .A2(
        interface3_bank_bus_dat_r[2]), .A3(interface4_bank_bus_dat_r[2]), .A4(
        interface6_bank_bus_dat_r[2]), .ZN(n715) );
  aoi22d1 U1341 ( .A1(n5394), .A2(mprj_dat_i[2]), .B1(n5395), .B2(
        mgmtsoc_vexriscv_debug_bus_dat_r[2]), .ZN(n714) );
  aon211d1 U1342 ( .C1(n716), .C2(n715), .B(n5356), .A(n714), .ZN(n717) );
  inv0d0 U1343 ( .I(n717), .ZN(n719) );
  buffd1 U1344 ( .I(n5380), .Z(n5437) );
  aoi22d1 U1345 ( .A1(n5437), .A2(\RAM256/Do0_pre[1][2] ), .B1(n5435), .B2(
        \RAM256/Do0_pre[0][2] ), .ZN(n718) );
  nd02d0 U1346 ( .A1(mprj_adr_o[5]), .A2(n722), .ZN(n728) );
  nr02d1 U1347 ( .A1(n725), .A2(n728), .ZN(n935) );
  nr02d1 U1348 ( .A1(n728), .A2(n1786), .ZN(n971) );
  aoi22d1 U1349 ( .A1(n935), .A2(n54), .B1(n971), .B2(n118), .ZN(n736) );
  inv0d0 U1350 ( .I(n2372), .ZN(n2373) );
  nr02d1 U1351 ( .A1(n727), .A2(n729), .ZN(n890) );
  nr02d1 U1352 ( .A1(n2451), .A2(n729), .ZN(n966) );
  aoi22d1 U1353 ( .A1(n890), .A2(csrbank6_oe1_w[16]), .B1(n966), .B2(
        csrbank6_ien0_w[16]), .ZN(n735) );
  nr02d0 U1354 ( .A1(mprj_adr_o[4]), .A2(n1783), .ZN(n1765) );
  buffd1 U1355 ( .I(n832), .Z(n936) );
  aoi22d1 U1356 ( .A1(n937), .A2(csrbank6_ien3_w[16]), .B1(n936), .B2(
        csrbank6_ien1_w[16]), .ZN(n734) );
  buffd1 U1357 ( .I(n737), .Z(n946) );
  inv0d0 U1358 ( .I(mprj_adr_o[5]), .ZN(n5621) );
  buffd1 U1359 ( .I(n945), .Z(n957) );
  aoi22d1 U1360 ( .A1(n946), .A2(csrbank6_oe3_w[16]), .B1(n957), .B2(n22), 
        .ZN(n732) );
  buffd1 U1361 ( .I(n875), .Z(n927) );
  aoi22d1 U1362 ( .A1(n919), .A2(csrbank6_oe2_w[16]), .B1(n927), .B2(
        csrbank6_ien2_w[16]), .ZN(n731) );
  buffd1 U1363 ( .I(n824), .Z(n2148) );
  aoi22d1 U1364 ( .A1(n947), .A2(n86), .B1(n2148), .B2(csrbank6_oe0_w[16]), 
        .ZN(n730) );
  an03d0 U1365 ( .A1(n732), .A2(n731), .A3(n730), .Z(n733) );
  aoi22d1 U1366 ( .A1(n947), .A2(n71), .B1(n971), .B2(n103), .ZN(n744) );
  buffd1 U1367 ( .I(n875), .Z(n970) );
  aoi22d1 U1368 ( .A1(n970), .A2(csrbank6_ien2_w[31]), .B1(n966), .B2(
        csrbank6_ien0_w[31]), .ZN(n743) );
  aoi22d1 U1369 ( .A1(n919), .A2(csrbank6_oe2_w[31]), .B1(n890), .B2(
        csrbank6_oe1_w[31]), .ZN(n742) );
  buffd1 U1370 ( .I(n935), .Z(n2067) );
  buffd1 U1371 ( .I(n737), .Z(n965) );
  aoi22d1 U1372 ( .A1(n2067), .A2(n39), .B1(n965), .B2(csrbank6_oe3_w[31]), 
        .ZN(n740) );
  buffd1 U1373 ( .I(n937), .Z(n2410) );
  buffd1 U1374 ( .I(n832), .Z(n969) );
  aoi22d1 U1375 ( .A1(n2410), .A2(csrbank6_ien3_w[31]), .B1(n969), .B2(
        csrbank6_ien1_w[31]), .ZN(n739) );
  aoi22d1 U1376 ( .A1(n957), .A2(n7), .B1(n2148), .B2(csrbank6_oe0_w[31]), 
        .ZN(n738) );
  an03d0 U1377 ( .A1(n740), .A2(n739), .A3(n738), .Z(n741) );
  buffd1 U1378 ( .I(n947), .Z(n2026) );
  aoi22d1 U1379 ( .A1(n935), .A2(n45), .B1(n2026), .B2(n77), .ZN(n753) );
  buffd1 U1380 ( .I(n919), .Z(n2221) );
  buffd1 U1381 ( .I(n937), .Z(n968) );
  aoi22d1 U1382 ( .A1(n2221), .A2(csrbank6_oe2_w[25]), .B1(n968), .B2(
        csrbank6_ien3_w[25]), .ZN(n752) );
  aoi22d1 U1383 ( .A1(n970), .A2(csrbank6_ien2_w[25]), .B1(n890), .B2(
        csrbank6_oe1_w[25]), .ZN(n751) );
  aoi22d1 U1384 ( .A1(n946), .A2(csrbank6_oe3_w[25]), .B1(n957), .B2(n13), 
        .ZN(n749) );
  aoi22d1 U1385 ( .A1(n966), .A2(csrbank6_ien0_w[25]), .B1(n969), .B2(
        csrbank6_ien1_w[25]), .ZN(n748) );
  buffd1 U1386 ( .I(n824), .Z(n967) );
  buffd1 U1387 ( .I(n971), .Z(n1985) );
  aoi22d1 U1388 ( .A1(n967), .A2(csrbank6_oe0_w[25]), .B1(n1985), .B2(n109), 
        .ZN(n747) );
  an03d0 U1389 ( .A1(n749), .A2(n748), .A3(n747), .Z(n750) );
  buffd3 U1390 ( .I(n1845), .Z(n4723) );
  inv0d0 U1391 ( .I(mgmtsoc_master_rxtx_w[29]), .ZN(n4716) );
  inv0d0 U1392 ( .I(mgmtsoc_master_rxtx_w[31]), .ZN(n4720) );
  nr02d0 U1393 ( .A1(n4723), .A2(n4720), .ZN(N4274) );
  inv0d0 U1394 ( .I(mgmtsoc_master_rxtx_w[30]), .ZN(n4719) );
  nr02d0 U1395 ( .A1(n4723), .A2(n4719), .ZN(N4273) );
  inv0d0 U1396 ( .I(mgmtsoc_master_rxtx_w[27]), .ZN(n4714) );
  nr02d0 U1397 ( .A1(n4723), .A2(n4714), .ZN(N4270) );
  inv0d0 U1398 ( .I(mgmtsoc_master_rxtx_w[26]), .ZN(n4713) );
  nr02d0 U1399 ( .A1(n4723), .A2(n4713), .ZN(N4269) );
  inv0d0 U1400 ( .I(mgmtsoc_master_rxtx_w[28]), .ZN(n4715) );
  inv0d0 U1401 ( .I(mgmtsoc_master_rxtx_w[25]), .ZN(n4712) );
  nr02d0 U1402 ( .A1(n4723), .A2(n4712), .ZN(N4268) );
  buffd1 U1403 ( .I(n947), .Z(n956) );
  aoi22d1 U1404 ( .A1(n957), .A2(n21), .B1(n956), .B2(n85), .ZN(n760) );
  aoi22d1 U1405 ( .A1(n890), .A2(csrbank6_oe1_w[17]), .B1(n966), .B2(
        csrbank6_ien0_w[17]), .ZN(n759) );
  aoi22d1 U1406 ( .A1(n2148), .A2(csrbank6_oe0_w[17]), .B1(n968), .B2(
        csrbank6_ien3_w[17]), .ZN(n758) );
  aoi22d1 U1407 ( .A1(n2067), .A2(n53), .B1(n965), .B2(csrbank6_oe3_w[17]), 
        .ZN(n756) );
  aoi22d1 U1408 ( .A1(n970), .A2(csrbank6_ien2_w[17]), .B1(n936), .B2(
        csrbank6_ien1_w[17]), .ZN(n755) );
  buffd1 U1409 ( .I(n919), .Z(n955) );
  aoi22d1 U1410 ( .A1(n955), .A2(csrbank6_oe2_w[17]), .B1(n1985), .B2(n117), 
        .ZN(n754) );
  an03d0 U1411 ( .A1(n756), .A2(n755), .A3(n754), .Z(n757) );
  aoi22d1 U1412 ( .A1(n945), .A2(n27), .B1(n956), .B2(n91), .ZN(n767) );
  aoi22d1 U1413 ( .A1(n970), .A2(csrbank6_ien2_w[11]), .B1(n966), .B2(
        csrbank6_ien0_w[11]), .ZN(n766) );
  aoi22d1 U1414 ( .A1(n890), .A2(csrbank6_oe1_w[11]), .B1(n936), .B2(
        csrbank6_ien1_w[11]), .ZN(n765) );
  aoi22d1 U1415 ( .A1(n935), .A2(n59), .B1(n965), .B2(csrbank6_oe3_w[11]), 
        .ZN(n763) );
  aoi22d1 U1416 ( .A1(n967), .A2(csrbank6_oe0_w[11]), .B1(n2410), .B2(
        csrbank6_ien3_w[11]), .ZN(n762) );
  aoi22d1 U1417 ( .A1(n955), .A2(csrbank6_oe2_w[11]), .B1(n1985), .B2(n123), 
        .ZN(n761) );
  an03d0 U1418 ( .A1(n763), .A2(n762), .A3(n761), .Z(n764) );
  aoi22d1 U1419 ( .A1(n935), .A2(n51), .B1(n945), .B2(n19), .ZN(n774) );
  aoi22d1 U1420 ( .A1(n970), .A2(csrbank6_ien2_w[19]), .B1(n966), .B2(
        csrbank6_ien0_w[19]), .ZN(n773) );
  aoi22d1 U1421 ( .A1(n890), .A2(csrbank6_oe1_w[19]), .B1(n969), .B2(
        csrbank6_ien1_w[19]), .ZN(n772) );
  aoi22d1 U1422 ( .A1(n965), .A2(csrbank6_oe3_w[19]), .B1(n956), .B2(n83), 
        .ZN(n770) );
  aoi22d1 U1423 ( .A1(n967), .A2(csrbank6_oe0_w[19]), .B1(n955), .B2(
        csrbank6_oe2_w[19]), .ZN(n769) );
  aoi22d1 U1424 ( .A1(n968), .A2(csrbank6_ien3_w[19]), .B1(n1985), .B2(n115), 
        .ZN(n768) );
  an03d0 U1425 ( .A1(n770), .A2(n769), .A3(n768), .Z(n771) );
  aoi22d1 U1426 ( .A1(n2067), .A2(n40), .B1(n2026), .B2(n72), .ZN(n781) );
  aoi22d1 U1427 ( .A1(n966), .A2(csrbank6_ien0_w[30]), .B1(n969), .B2(
        csrbank6_ien1_w[30]), .ZN(n780) );
  aoi22d1 U1428 ( .A1(n967), .A2(csrbank6_oe0_w[30]), .B1(n970), .B2(
        csrbank6_ien2_w[30]), .ZN(n779) );
  aoi22d1 U1429 ( .A1(n946), .A2(csrbank6_oe3_w[30]), .B1(n1985), .B2(n104), 
        .ZN(n777) );
  aoi22d1 U1430 ( .A1(n955), .A2(csrbank6_oe2_w[30]), .B1(n890), .B2(
        csrbank6_oe1_w[30]), .ZN(n776) );
  aoi22d1 U1431 ( .A1(n957), .A2(n8), .B1(n968), .B2(csrbank6_ien3_w[30]), 
        .ZN(n775) );
  an03d0 U1432 ( .A1(n777), .A2(n776), .A3(n775), .Z(n778) );
  buffd1 U1433 ( .I(n945), .Z(n2108) );
  aoi22d1 U1434 ( .A1(n946), .A2(csrbank6_oe3_w[24]), .B1(n2108), .B2(n14), 
        .ZN(n788) );
  aoi22d1 U1435 ( .A1(n967), .A2(csrbank6_oe0_w[24]), .B1(n890), .B2(
        csrbank6_oe1_w[24]), .ZN(n787) );
  aoi22d1 U1436 ( .A1(n966), .A2(csrbank6_ien0_w[24]), .B1(n969), .B2(
        csrbank6_ien1_w[24]), .ZN(n786) );
  aoi22d1 U1437 ( .A1(n935), .A2(n46), .B1(n971), .B2(n110), .ZN(n784) );
  aoi22d1 U1438 ( .A1(n955), .A2(csrbank6_oe2_w[24]), .B1(n927), .B2(
        csrbank6_ien2_w[24]), .ZN(n783) );
  aoi22d1 U1439 ( .A1(n947), .A2(n78), .B1(n968), .B2(csrbank6_ien3_w[24]), 
        .ZN(n782) );
  an03d0 U1440 ( .A1(n784), .A2(n783), .A3(n782), .Z(n785) );
  aoi22d1 U1441 ( .A1(n935), .A2(n68), .B1(n1985), .B2(n132), .ZN(n795) );
  aoi22d1 U1442 ( .A1(n2148), .A2(csrbank6_oe0_w[2]), .B1(n937), .B2(
        csrbank6_ien3_w[2]), .ZN(n794) );
  buffd1 U1443 ( .I(n890), .Z(n2183) );
  aoi22d1 U1444 ( .A1(n2183), .A2(csrbank6_oe1_w[2]), .B1(n966), .B2(
        csrbank6_ien0_w[2]), .ZN(n793) );
  aoi22d1 U1445 ( .A1(n946), .A2(csrbank6_oe3_w[2]), .B1(n957), .B2(n36), .ZN(
        n791) );
  aoi22d1 U1446 ( .A1(n927), .A2(csrbank6_ien2_w[2]), .B1(n936), .B2(
        csrbank6_ien1_w[2]), .ZN(n790) );
  aoi22d1 U1447 ( .A1(n956), .A2(n100), .B1(n2221), .B2(csrbank6_oe2_w[2]), 
        .ZN(n789) );
  an03d0 U1448 ( .A1(n791), .A2(n790), .A3(n789), .Z(n792) );
  aoi22d1 U1449 ( .A1(n946), .A2(csrbank6_oe3_w[13]), .B1(n2108), .B2(n25), 
        .ZN(n802) );
  aoi22d1 U1450 ( .A1(n968), .A2(csrbank6_ien3_w[13]), .B1(n2183), .B2(
        csrbank6_oe1_w[13]), .ZN(n801) );
  aoi22d1 U1451 ( .A1(n966), .A2(csrbank6_ien0_w[13]), .B1(n936), .B2(
        csrbank6_ien1_w[13]), .ZN(n800) );
  aoi22d1 U1452 ( .A1(n935), .A2(n57), .B1(n1985), .B2(n121), .ZN(n798) );
  aoi22d1 U1453 ( .A1(n967), .A2(csrbank6_oe0_w[13]), .B1(n955), .B2(
        csrbank6_oe2_w[13]), .ZN(n797) );
  aoi22d1 U1454 ( .A1(n2026), .A2(n89), .B1(n927), .B2(csrbank6_ien2_w[13]), 
        .ZN(n796) );
  an03d0 U1455 ( .A1(n798), .A2(n797), .A3(n796), .Z(n799) );
  aoi22d1 U1456 ( .A1(n946), .A2(csrbank6_oe3_w[15]), .B1(n971), .B2(n119), 
        .ZN(n809) );
  aoi22d1 U1457 ( .A1(n970), .A2(csrbank6_ien2_w[15]), .B1(n2183), .B2(
        csrbank6_oe1_w[15]), .ZN(n808) );
  aoi22d1 U1458 ( .A1(n966), .A2(csrbank6_ien0_w[15]), .B1(n936), .B2(
        csrbank6_ien1_w[15]), .ZN(n807) );
  aoi22d1 U1459 ( .A1(n2108), .A2(n23), .B1(n956), .B2(n87), .ZN(n805) );
  aoi22d1 U1460 ( .A1(n967), .A2(csrbank6_oe0_w[15]), .B1(n968), .B2(
        csrbank6_ien3_w[15]), .ZN(n804) );
  aoi22d1 U1461 ( .A1(n2067), .A2(n55), .B1(n955), .B2(csrbank6_oe2_w[15]), 
        .ZN(n803) );
  an03d0 U1462 ( .A1(n805), .A2(n804), .A3(n803), .Z(n806) );
  aoi22d1 U1463 ( .A1(n946), .A2(csrbank6_oe3_w[5]), .B1(n2108), .B2(n33), 
        .ZN(n816) );
  buffd1 U1464 ( .I(n966), .Z(n2295) );
  aoi22d1 U1465 ( .A1(n2148), .A2(csrbank6_oe0_w[5]), .B1(n2295), .B2(
        csrbank6_ien0_w[5]), .ZN(n815) );
  aoi22d1 U1466 ( .A1(n890), .A2(csrbank6_oe1_w[5]), .B1(n969), .B2(
        csrbank6_ien1_w[5]), .ZN(n814) );
  aoi22d1 U1467 ( .A1(n956), .A2(n97), .B1(n1985), .B2(n129), .ZN(n812) );
  aoi22d1 U1468 ( .A1(n955), .A2(csrbank6_oe2_w[5]), .B1(n2410), .B2(
        csrbank6_ien3_w[5]), .ZN(n811) );
  aoi22d1 U1469 ( .A1(n2067), .A2(n65), .B1(n927), .B2(csrbank6_ien2_w[5]), 
        .ZN(n810) );
  an03d0 U1470 ( .A1(n812), .A2(n811), .A3(n810), .Z(n813) );
  aoi22d1 U1471 ( .A1(n956), .A2(n98), .B1(n1985), .B2(n130), .ZN(n823) );
  aoi22d1 U1472 ( .A1(n967), .A2(csrbank6_oe0_w[4]), .B1(n2221), .B2(
        csrbank6_oe2_w[4]), .ZN(n822) );
  aoi22d1 U1473 ( .A1(n2410), .A2(csrbank6_ien3_w[4]), .B1(n2295), .B2(
        csrbank6_ien0_w[4]), .ZN(n821) );
  aoi22d1 U1474 ( .A1(n2067), .A2(n66), .B1(n2108), .B2(n34), .ZN(n819) );
  aoi22d1 U1475 ( .A1(n890), .A2(csrbank6_oe1_w[4]), .B1(n936), .B2(
        csrbank6_ien1_w[4]), .ZN(n818) );
  aoi22d1 U1476 ( .A1(n946), .A2(csrbank6_oe3_w[4]), .B1(n927), .B2(
        csrbank6_ien2_w[4]), .ZN(n817) );
  an03d0 U1477 ( .A1(n819), .A2(n818), .A3(n817), .Z(n820) );
  aoi22d1 U1478 ( .A1(n965), .A2(csrbank6_oe3_w[21]), .B1(n945), .B2(n17), 
        .ZN(n831) );
  aoi22d1 U1479 ( .A1(n890), .A2(csrbank6_oe1_w[21]), .B1(n936), .B2(
        csrbank6_ien1_w[21]), .ZN(n830) );
  aoi22d1 U1480 ( .A1(n824), .A2(csrbank6_oe0_w[21]), .B1(n2295), .B2(
        csrbank6_ien0_w[21]), .ZN(n829) );
  aoi22d1 U1481 ( .A1(n935), .A2(n49), .B1(n1985), .B2(n113), .ZN(n827) );
  aoi22d1 U1482 ( .A1(n968), .A2(csrbank6_ien3_w[21]), .B1(n970), .B2(
        csrbank6_ien2_w[21]), .ZN(n826) );
  aoi22d1 U1483 ( .A1(n947), .A2(n81), .B1(n955), .B2(csrbank6_oe2_w[21]), 
        .ZN(n825) );
  an03d0 U1484 ( .A1(n827), .A2(n826), .A3(n825), .Z(n828) );
  aoi22d1 U1485 ( .A1(n965), .A2(csrbank6_oe3_w[22]), .B1(n945), .B2(n16), 
        .ZN(n839) );
  aoi22d1 U1486 ( .A1(n927), .A2(csrbank6_ien2_w[22]), .B1(n832), .B2(
        csrbank6_ien1_w[22]), .ZN(n838) );
  aoi22d1 U1487 ( .A1(n955), .A2(csrbank6_oe2_w[22]), .B1(n2295), .B2(
        csrbank6_ien0_w[22]), .ZN(n837) );
  aoi22d1 U1488 ( .A1(n935), .A2(n48), .B1(n1985), .B2(n112), .ZN(n835) );
  aoi22d1 U1489 ( .A1(n967), .A2(csrbank6_oe0_w[22]), .B1(n890), .B2(
        csrbank6_oe1_w[22]), .ZN(n834) );
  aoi22d1 U1490 ( .A1(n947), .A2(n80), .B1(n968), .B2(csrbank6_ien3_w[22]), 
        .ZN(n833) );
  an03d0 U1491 ( .A1(n835), .A2(n834), .A3(n833), .Z(n836) );
  aoi22d1 U1492 ( .A1(n957), .A2(n11), .B1(n2026), .B2(n75), .ZN(n846) );
  aoi22d1 U1493 ( .A1(n2410), .A2(csrbank6_ien3_w[27]), .B1(n890), .B2(
        csrbank6_oe1_w[27]), .ZN(n845) );
  aoi22d1 U1494 ( .A1(n919), .A2(csrbank6_oe2_w[27]), .B1(n2295), .B2(
        csrbank6_ien0_w[27]), .ZN(n844) );
  aoi22d1 U1495 ( .A1(n2067), .A2(n43), .B1(n965), .B2(csrbank6_oe3_w[27]), 
        .ZN(n842) );
  aoi22d1 U1496 ( .A1(n967), .A2(csrbank6_oe0_w[27]), .B1(n970), .B2(
        csrbank6_ien2_w[27]), .ZN(n841) );
  aoi22d1 U1497 ( .A1(n971), .A2(n107), .B1(n969), .B2(csrbank6_ien1_w[27]), 
        .ZN(n840) );
  an03d0 U1498 ( .A1(n842), .A2(n841), .A3(n840), .Z(n843) );
  aoi22d1 U1499 ( .A1(n935), .A2(n67), .B1(n965), .B2(csrbank6_oe3_w[3]), .ZN(
        n853) );
  aoi22d1 U1500 ( .A1(n2148), .A2(csrbank6_oe0_w[3]), .B1(n2410), .B2(
        csrbank6_ien3_w[3]), .ZN(n852) );
  aoi22d1 U1501 ( .A1(n919), .A2(csrbank6_oe2_w[3]), .B1(n2183), .B2(
        csrbank6_oe1_w[3]), .ZN(n851) );
  aoi22d1 U1502 ( .A1(n957), .A2(n35), .B1(n1985), .B2(n131), .ZN(n849) );
  aoi22d1 U1503 ( .A1(n966), .A2(csrbank6_ien0_w[3]), .B1(n969), .B2(
        csrbank6_ien1_w[3]), .ZN(n848) );
  aoi22d1 U1504 ( .A1(n956), .A2(n99), .B1(n927), .B2(csrbank6_ien2_w[3]), 
        .ZN(n847) );
  an03d0 U1505 ( .A1(n849), .A2(n848), .A3(n847), .Z(n850) );
  aoi22d1 U1506 ( .A1(n957), .A2(n37), .B1(n971), .B2(n133), .ZN(n860) );
  aoi22d1 U1507 ( .A1(n2295), .A2(csrbank6_ien0_w[1]), .B1(n936), .B2(
        csrbank6_ien1_w[1]), .ZN(n859) );
  aoi22d1 U1508 ( .A1(n937), .A2(csrbank6_ien3_w[1]), .B1(n2183), .B2(
        csrbank6_oe1_w[1]), .ZN(n858) );
  aoi22d1 U1509 ( .A1(n946), .A2(csrbank6_oe3_w[1]), .B1(n2026), .B2(n101), 
        .ZN(n856) );
  aoi22d1 U1510 ( .A1(n2148), .A2(csrbank6_oe0_w[1]), .B1(n2221), .B2(
        csrbank6_oe2_w[1]), .ZN(n855) );
  aoi22d1 U1511 ( .A1(n2067), .A2(n69), .B1(n970), .B2(csrbank6_ien2_w[1]), 
        .ZN(n854) );
  an03d0 U1512 ( .A1(n856), .A2(n855), .A3(n854), .Z(n857) );
  aoi22d1 U1513 ( .A1(n957), .A2(n31), .B1(n1985), .B2(n127), .ZN(n867) );
  aoi22d1 U1514 ( .A1(n2148), .A2(csrbank6_oe0_w[7]), .B1(n2221), .B2(
        csrbank6_oe2_w[7]), .ZN(n866) );
  aoi22d1 U1515 ( .A1(n890), .A2(csrbank6_oe1_w[7]), .B1(n936), .B2(
        csrbank6_ien1_w[7]), .ZN(n865) );
  aoi22d1 U1516 ( .A1(n946), .A2(csrbank6_oe3_w[7]), .B1(n956), .B2(n95), .ZN(
        n863) );
  aoi22d1 U1517 ( .A1(n968), .A2(csrbank6_ien3_w[7]), .B1(n2295), .B2(
        csrbank6_ien0_w[7]), .ZN(n862) );
  aoi22d1 U1518 ( .A1(n935), .A2(n63), .B1(n927), .B2(csrbank6_ien2_w[7]), 
        .ZN(n861) );
  an03d0 U1519 ( .A1(n863), .A2(n862), .A3(n861), .Z(n864) );
  aoi22d1 U1520 ( .A1(n935), .A2(n44), .B1(n971), .B2(n108), .ZN(n874) );
  aoi22d1 U1521 ( .A1(n970), .A2(csrbank6_ien2_w[26]), .B1(n966), .B2(
        csrbank6_ien0_w[26]), .ZN(n873) );
  aoi22d1 U1522 ( .A1(n919), .A2(csrbank6_oe2_w[26]), .B1(n968), .B2(
        csrbank6_ien3_w[26]), .ZN(n872) );
  aoi22d1 U1523 ( .A1(n957), .A2(n12), .B1(n956), .B2(n76), .ZN(n870) );
  aoi22d1 U1524 ( .A1(n967), .A2(csrbank6_oe0_w[26]), .B1(n2183), .B2(
        csrbank6_oe1_w[26]), .ZN(n869) );
  aoi22d1 U1525 ( .A1(n946), .A2(csrbank6_oe3_w[26]), .B1(n969), .B2(
        csrbank6_ien1_w[26]), .ZN(n868) );
  an03d0 U1526 ( .A1(n870), .A2(n869), .A3(n868), .Z(n871) );
  aoi22d1 U1527 ( .A1(n946), .A2(csrbank6_oe3_w[20]), .B1(n2026), .B2(n82), 
        .ZN(n882) );
  aoi22d1 U1528 ( .A1(n2148), .A2(csrbank6_oe0_w[20]), .B1(n890), .B2(
        csrbank6_oe1_w[20]), .ZN(n881) );
  aoi22d1 U1529 ( .A1(n875), .A2(csrbank6_ien2_w[20]), .B1(n936), .B2(
        csrbank6_ien1_w[20]), .ZN(n880) );
  aoi22d1 U1530 ( .A1(n957), .A2(n18), .B1(n971), .B2(n114), .ZN(n878) );
  aoi22d1 U1531 ( .A1(n955), .A2(csrbank6_oe2_w[20]), .B1(n2295), .B2(
        csrbank6_ien0_w[20]), .ZN(n877) );
  aoi22d1 U1532 ( .A1(n2067), .A2(n50), .B1(n968), .B2(csrbank6_ien3_w[20]), 
        .ZN(n876) );
  an03d0 U1533 ( .A1(n878), .A2(n877), .A3(n876), .Z(n879) );
  aoi22d1 U1534 ( .A1(n957), .A2(n15), .B1(n1985), .B2(n111), .ZN(n889) );
  aoi22d1 U1535 ( .A1(n955), .A2(csrbank6_oe2_w[23]), .B1(n2295), .B2(
        csrbank6_ien0_w[23]), .ZN(n888) );
  aoi22d1 U1536 ( .A1(n937), .A2(csrbank6_ien3_w[23]), .B1(n969), .B2(
        csrbank6_ien1_w[23]), .ZN(n887) );
  aoi22d1 U1537 ( .A1(n965), .A2(csrbank6_oe3_w[23]), .B1(n956), .B2(n79), 
        .ZN(n885) );
  aoi22d1 U1538 ( .A1(n967), .A2(csrbank6_oe0_w[23]), .B1(n2183), .B2(
        csrbank6_oe1_w[23]), .ZN(n884) );
  aoi22d1 U1539 ( .A1(n2067), .A2(n47), .B1(n927), .B2(csrbank6_ien2_w[23]), 
        .ZN(n883) );
  an03d0 U1540 ( .A1(n885), .A2(n884), .A3(n883), .Z(n886) );
  aoi22d1 U1541 ( .A1(n935), .A2(n56), .B1(n2108), .B2(n24), .ZN(n897) );
  aoi22d1 U1542 ( .A1(n2148), .A2(csrbank6_oe0_w[14]), .B1(n890), .B2(
        csrbank6_oe1_w[14]), .ZN(n896) );
  aoi22d1 U1543 ( .A1(n2410), .A2(csrbank6_ien3_w[14]), .B1(n927), .B2(
        csrbank6_ien2_w[14]), .ZN(n895) );
  aoi22d1 U1544 ( .A1(n965), .A2(csrbank6_oe3_w[14]), .B1(n956), .B2(n88), 
        .ZN(n893) );
  aoi22d1 U1545 ( .A1(n2221), .A2(csrbank6_oe2_w[14]), .B1(n2295), .B2(
        csrbank6_ien0_w[14]), .ZN(n892) );
  aoi22d1 U1546 ( .A1(n971), .A2(n120), .B1(n936), .B2(csrbank6_ien1_w[14]), 
        .ZN(n891) );
  an03d0 U1547 ( .A1(n893), .A2(n892), .A3(n891), .Z(n894) );
  aoi22d1 U1548 ( .A1(n935), .A2(n62), .B1(n946), .B2(csrbank6_oe3_w[8]), .ZN(
        n904) );
  aoi22d1 U1549 ( .A1(n2148), .A2(csrbank6_oe0_w[8]), .B1(n955), .B2(
        csrbank6_oe2_w[8]), .ZN(n903) );
  aoi22d1 U1550 ( .A1(n966), .A2(csrbank6_ien0_w[8]), .B1(n969), .B2(
        csrbank6_ien1_w[8]), .ZN(n902) );
  aoi22d1 U1551 ( .A1(n957), .A2(n30), .B1(n971), .B2(n126), .ZN(n900) );
  aoi22d1 U1552 ( .A1(n968), .A2(csrbank6_ien3_w[8]), .B1(n2183), .B2(
        csrbank6_oe1_w[8]), .ZN(n899) );
  aoi22d1 U1553 ( .A1(n956), .A2(n94), .B1(n927), .B2(csrbank6_ien2_w[8]), 
        .ZN(n898) );
  an03d0 U1554 ( .A1(n900), .A2(n899), .A3(n898), .Z(n901) );
  aoi22d1 U1555 ( .A1(n957), .A2(n32), .B1(n971), .B2(n128), .ZN(n911) );
  aoi22d1 U1556 ( .A1(n967), .A2(csrbank6_oe0_w[6]), .B1(n969), .B2(
        csrbank6_ien1_w[6]), .ZN(n910) );
  aoi22d1 U1557 ( .A1(n968), .A2(csrbank6_ien3_w[6]), .B1(n2295), .B2(
        csrbank6_ien0_w[6]), .ZN(n909) );
  aoi22d1 U1558 ( .A1(n2067), .A2(n64), .B1(n965), .B2(csrbank6_oe3_w[6]), 
        .ZN(n907) );
  aoi22d1 U1559 ( .A1(n927), .A2(csrbank6_ien2_w[6]), .B1(n2183), .B2(
        csrbank6_oe1_w[6]), .ZN(n906) );
  aoi22d1 U1560 ( .A1(n956), .A2(n96), .B1(n2221), .B2(csrbank6_oe2_w[6]), 
        .ZN(n905) );
  an03d0 U1561 ( .A1(n907), .A2(n906), .A3(n905), .Z(n908) );
  aoi22d1 U1562 ( .A1(n2108), .A2(n28), .B1(n971), .B2(n124), .ZN(n918) );
  aoi22d1 U1563 ( .A1(n937), .A2(csrbank6_ien3_w[10]), .B1(n2183), .B2(
        csrbank6_oe1_w[10]), .ZN(n917) );
  aoi22d1 U1564 ( .A1(n2148), .A2(csrbank6_oe0_w[10]), .B1(n970), .B2(
        csrbank6_ien2_w[10]), .ZN(n916) );
  aoi22d1 U1565 ( .A1(n965), .A2(csrbank6_oe3_w[10]), .B1(n956), .B2(n92), 
        .ZN(n914) );
  aoi22d1 U1566 ( .A1(n2221), .A2(csrbank6_oe2_w[10]), .B1(n2295), .B2(
        csrbank6_ien0_w[10]), .ZN(n913) );
  aoi22d1 U1567 ( .A1(n2067), .A2(n60), .B1(n936), .B2(csrbank6_ien1_w[10]), 
        .ZN(n912) );
  an03d0 U1568 ( .A1(n914), .A2(n913), .A3(n912), .Z(n915) );
  aoi22d1 U1569 ( .A1(n2026), .A2(n90), .B1(n971), .B2(n122), .ZN(n926) );
  aoi22d1 U1570 ( .A1(n2148), .A2(csrbank6_oe0_w[12]), .B1(n927), .B2(
        csrbank6_ien2_w[12]), .ZN(n925) );
  aoi22d1 U1571 ( .A1(n919), .A2(csrbank6_oe2_w[12]), .B1(n936), .B2(
        csrbank6_ien1_w[12]), .ZN(n924) );
  aoi22d1 U1572 ( .A1(n965), .A2(csrbank6_oe3_w[12]), .B1(n2108), .B2(n26), 
        .ZN(n922) );
  aoi22d1 U1573 ( .A1(n2183), .A2(csrbank6_oe1_w[12]), .B1(n2295), .B2(
        csrbank6_ien0_w[12]), .ZN(n921) );
  aoi22d1 U1574 ( .A1(n2067), .A2(n58), .B1(n2410), .B2(csrbank6_ien3_w[12]), 
        .ZN(n920) );
  aoi22d1 U1575 ( .A1(n935), .A2(n61), .B1(n2108), .B2(n29), .ZN(n934) );
  aoi22d1 U1576 ( .A1(n955), .A2(csrbank6_oe2_w[9]), .B1(n2410), .B2(
        csrbank6_ien3_w[9]), .ZN(n933) );
  aoi22d1 U1577 ( .A1(n967), .A2(csrbank6_oe0_w[9]), .B1(n927), .B2(
        csrbank6_ien2_w[9]), .ZN(n932) );
  aoi22d1 U1578 ( .A1(n946), .A2(csrbank6_oe3_w[9]), .B1(n956), .B2(n93), .ZN(
        n930) );
  aoi22d1 U1579 ( .A1(n2183), .A2(csrbank6_oe1_w[9]), .B1(n2295), .B2(
        csrbank6_ien0_w[9]), .ZN(n929) );
  aoi22d1 U1580 ( .A1(n971), .A2(n125), .B1(n936), .B2(csrbank6_ien1_w[9]), 
        .ZN(n928) );
  aoi22d1 U1581 ( .A1(n935), .A2(n52), .B1(n965), .B2(csrbank6_oe3_w[18]), 
        .ZN(n944) );
  aoi22d1 U1582 ( .A1(n2148), .A2(csrbank6_oe0_w[18]), .B1(n955), .B2(
        csrbank6_oe2_w[18]), .ZN(n943) );
  aoi22d1 U1583 ( .A1(n937), .A2(csrbank6_ien3_w[18]), .B1(n936), .B2(
        csrbank6_ien1_w[18]), .ZN(n942) );
  aoi22d1 U1584 ( .A1(n957), .A2(n20), .B1(n1985), .B2(n116), .ZN(n940) );
  aoi22d1 U1585 ( .A1(n970), .A2(csrbank6_ien2_w[18]), .B1(n2295), .B2(
        csrbank6_ien0_w[18]), .ZN(n939) );
  aoi22d1 U1586 ( .A1(n2026), .A2(n84), .B1(n2183), .B2(csrbank6_oe1_w[18]), 
        .ZN(n938) );
  an03d0 U1587 ( .A1(n940), .A2(n939), .A3(n938), .Z(n941) );
  aoi22d1 U1588 ( .A1(n946), .A2(csrbank6_oe3_w[29]), .B1(n945), .B2(n9), .ZN(
        n954) );
  aoi22d1 U1589 ( .A1(n967), .A2(csrbank6_oe0_w[29]), .B1(n955), .B2(
        csrbank6_oe2_w[29]), .ZN(n953) );
  aoi22d1 U1590 ( .A1(n966), .A2(csrbank6_ien0_w[29]), .B1(n969), .B2(
        csrbank6_ien1_w[29]), .ZN(n952) );
  aoi22d1 U1591 ( .A1(n947), .A2(n73), .B1(n1985), .B2(n105), .ZN(n950) );
  aoi22d1 U1592 ( .A1(n968), .A2(csrbank6_ien3_w[29]), .B1(n970), .B2(
        csrbank6_ien2_w[29]), .ZN(n949) );
  aoi22d1 U1593 ( .A1(n2067), .A2(n41), .B1(n2183), .B2(csrbank6_oe1_w[29]), 
        .ZN(n948) );
  an03d0 U1594 ( .A1(n950), .A2(n949), .A3(n948), .Z(n951) );
  aoi22d1 U1595 ( .A1(n2067), .A2(n70), .B1(csrbank6_oe3_w[0]), .B2(n965), 
        .ZN(n964) );
  aoi22d1 U1596 ( .A1(n968), .A2(csrbank6_ien3_w[0]), .B1(csrbank6_ien2_w[0]), 
        .B2(n970), .ZN(n963) );
  aoi22d1 U1597 ( .A1(n967), .A2(csrbank6_oe0_w[0]), .B1(n955), .B2(
        csrbank6_oe2_w[0]), .ZN(n962) );
  aoi22d1 U1598 ( .A1(n957), .A2(n38), .B1(n956), .B2(n102), .ZN(n960) );
  aoi22d1 U1599 ( .A1(n2295), .A2(csrbank6_ien0_w[0]), .B1(csrbank6_ien1_w[0]), 
        .B2(n969), .ZN(n959) );
  aoi22d1 U1600 ( .A1(n971), .A2(n134), .B1(n2183), .B2(csrbank6_oe1_w[0]), 
        .ZN(n958) );
  an03d0 U1601 ( .A1(n960), .A2(n959), .A3(n958), .Z(n961) );
  aoi22d1 U1602 ( .A1(n2067), .A2(n42), .B1(n965), .B2(csrbank6_oe3_w[28]), 
        .ZN(n978) );
  aoi22d1 U1603 ( .A1(n967), .A2(csrbank6_oe0_w[28]), .B1(n966), .B2(
        csrbank6_ien0_w[28]), .ZN(n977) );
  aoi22d1 U1604 ( .A1(n2221), .A2(csrbank6_oe2_w[28]), .B1(n968), .B2(
        csrbank6_ien3_w[28]), .ZN(n976) );
  aoi22d1 U1605 ( .A1(n2108), .A2(n10), .B1(n2026), .B2(n74), .ZN(n974) );
  aoi22d1 U1606 ( .A1(n970), .A2(csrbank6_ien2_w[28]), .B1(n969), .B2(
        csrbank6_ien1_w[28]), .ZN(n973) );
  aoi22d1 U1607 ( .A1(n971), .A2(n106), .B1(n2183), .B2(csrbank6_oe1_w[28]), 
        .ZN(n972) );
  an03d0 U1608 ( .A1(n974), .A2(n973), .A3(n972), .Z(n975) );
  an02d0 U1609 ( .A1(n993), .A2(n980), .Z(N5446) );
  ah01d1 U1610 ( .A(n981), .B(mgmtsoc_litespisdrphycore_cnt[3]), .CO(n986), 
        .S(n980) );
  xr02d1 U1611 ( .A1(n982), .A2(mgmtsoc_litespisdrphycore_cnt[7]), .Z(n983) );
  an02d0 U1612 ( .A1(n993), .A2(n983), .Z(N5450) );
  ah01d1 U1613 ( .A(n984), .B(mgmtsoc_litespisdrphycore_cnt[5]), .CO(n991), 
        .S(n985) );
  an02d0 U1614 ( .A1(n993), .A2(n985), .Z(N5448) );
  ah01d1 U1615 ( .A(n986), .B(mgmtsoc_litespisdrphycore_cnt[4]), .CO(n984), 
        .S(n987) );
  an02d0 U1616 ( .A1(n993), .A2(n987), .Z(N5447) );
  ah01d1 U1617 ( .A(mgmtsoc_litespisdrphycore_cnt[0]), .B(
        mgmtsoc_litespisdrphycore_cnt[1]), .CO(n989), .S(n988) );
  an02d0 U1618 ( .A1(n993), .A2(n988), .Z(N5444) );
  ah01d1 U1619 ( .A(n989), .B(mgmtsoc_litespisdrphycore_cnt[2]), .CO(n981), 
        .S(n990) );
  an02d0 U1620 ( .A1(n993), .A2(n990), .Z(N5445) );
  ah01d1 U1621 ( .A(n991), .B(mgmtsoc_litespisdrphycore_cnt[6]), .CO(n982), 
        .S(n992) );
  an02d0 U1622 ( .A1(n993), .A2(n992), .Z(N5449) );
  an02d0 U1623 ( .A1(n2557), .A2(uart_rx_fifo_fifo_out_payload_data[3]), .Z(
        N4775) );
  an02d0 U1624 ( .A1(n2557), .A2(uart_rx_fifo_fifo_out_payload_data[2]), .Z(
        N4774) );
  an02d0 U1625 ( .A1(n2557), .A2(uart_rx_fifo_fifo_out_payload_data[4]), .Z(
        N4776) );
  an02d0 U1626 ( .A1(n2557), .A2(uart_rx_fifo_fifo_out_payload_data[5]), .Z(
        N4777) );
  an02d0 U1627 ( .A1(n2557), .A2(uart_rx_fifo_fifo_out_payload_data[7]), .Z(
        N4779) );
  an02d0 U1628 ( .A1(n2557), .A2(uart_rx_fifo_fifo_out_payload_data[6]), .Z(
        N4778) );
  inv0d0 U1629 ( .I(dbg_uart_dbg_uart_tx), .ZN(n2510) );
  aoim22d1 U1630 ( .A1(debug_in), .A2(n2510), .B1(sys_uart_tx), .B2(debug_in), 
        .Z(serial_tx) );
  an02d0 U1631 ( .A1(mgmtsoc_zero1), .A2(mgmtsoc_zero2), .Z(
        mgmtsoc_interrupt[0]) );
  an02d0 U1632 ( .A1(gpioin5_i02), .A2(gpioin5_i01), .Z(mgmtsoc_interrupt[7])
         );
  an02d0 U1633 ( .A1(gpioin3_i02), .A2(gpioin3_i01), .Z(mgmtsoc_interrupt[5])
         );
  an02d0 U1634 ( .A1(gpioin4_i02), .A2(gpioin4_i01), .Z(mgmtsoc_interrupt[6])
         );
  an02d0 U1635 ( .A1(gpioin2_i02), .A2(gpioin2_i01), .Z(mgmtsoc_interrupt[4])
         );
  an02d0 U1636 ( .A1(gpioin1_i01), .A2(gpioin1_i02), .Z(mgmtsoc_interrupt[3])
         );
  an02d0 U1637 ( .A1(gpioin0_i02), .A2(gpioin0_i01), .Z(mgmtsoc_interrupt[2])
         );
  ah01d1 U1638 ( .A(n994), .B(uart_phy_tx_phase[7]), .CO(n997), .S(n995) );
  an02d0 U1639 ( .A1(rs232phy_rs232phytx_state), .A2(n995), .Z(N3579) );
  ah01d1 U1640 ( .A(uart_phy_tx_phase[5]), .B(uart_phy_tx_phase[6]), .CO(n994), 
        .S(n996) );
  an02d0 U1641 ( .A1(rs232phy_rs232phytx_state), .A2(n996), .Z(N3578) );
  ah01d1 U1642 ( .A(n997), .B(uart_phy_tx_phase[8]), .CO(n1464), .S(n998) );
  an02d0 U1643 ( .A1(rs232phy_rs232phytx_state), .A2(n998), .Z(N3580) );
  inv0d0 U1644 ( .I(uart_phy_rx_phase[5]), .ZN(n999) );
  an02d0 U1645 ( .A1(rs232phy_rs232phyrx_state), .A2(n999), .Z(N3644) );
  ah01d1 U1646 ( .A(uart_phy_rx_phase[5]), .B(uart_phy_rx_phase[6]), .CO(n1001), .S(n1000) );
  an02d0 U1647 ( .A1(rs232phy_rs232phyrx_state), .A2(n1000), .Z(N3645) );
  ah01d1 U1648 ( .A(n1001), .B(uart_phy_rx_phase[7]), .CO(n1003), .S(n1002) );
  an02d0 U1649 ( .A1(rs232phy_rs232phyrx_state), .A2(n1002), .Z(N3646) );
  ah01d1 U1650 ( .A(n1003), .B(uart_phy_rx_phase[8]), .CO(n1006), .S(n1004) );
  an02d0 U1651 ( .A1(rs232phy_rs232phyrx_state), .A2(n1004), .Z(N3647) );
  aoi22d1 U1652 ( .A1(uart_phy_rx_phase[9]), .A2(n1007), .B1(n1006), .B2(n1005), .ZN(n1008) );
  an02d0 U1653 ( .A1(rs232phy_rs232phyrx_state), .A2(n1008), .Z(N3648) );
  an02d0 U1654 ( .A1(debug_in), .A2(serial_rx), .Z(dbg_uart_dbg_uart_rx) );
  or02d0 U1655 ( .A1(uart_enabled_o), .A2(debug_in), .Z(uart_enabled) );
  ah01d1 U1656 ( .A(n1009), .B(uart_phy_tx_phase[10]), .CO(n674), .S(n1010) );
  an02d0 U1657 ( .A1(rs232phy_rs232phytx_state), .A2(n1010), .Z(N3582) );
  aoi22d1 U1658 ( .A1(uart_phy_rx_phase[11]), .A2(n1013), .B1(n1012), .B2(
        n1011), .ZN(n1014) );
  an02d0 U1659 ( .A1(rs232phy_rs232phyrx_state), .A2(n1014), .Z(N3650) );
  ah01d1 U1660 ( .A(n1015), .B(uart_phy_rx_phase[10]), .CO(n1012), .S(n1016)
         );
  an02d0 U1661 ( .A1(n1200), .A2(n1016), .Z(N3649) );
  ah01d1 U1662 ( .A(n1017), .B(uart_phy_rx_phase[12]), .CO(n1022), .S(n1018)
         );
  an02d0 U1663 ( .A1(n1200), .A2(n1018), .Z(N3651) );
  inv0d0 U1664 ( .I(uart_phy_rx_phase[14]), .ZN(n1020) );
  nr02d0 U1665 ( .A1(uart_phy_rx_phase[13]), .A2(n1022), .ZN(n1019) );
  mx02d1 U1666 ( .I0(uart_phy_rx_phase[14]), .I1(n1020), .S(n1019), .Z(n1021)
         );
  an02d0 U1667 ( .A1(n1200), .A2(n1021), .Z(N3653) );
  inv0d0 U1668 ( .I(n1022), .ZN(n1023) );
  aoim22d1 U1669 ( .A1(uart_phy_rx_phase[13]), .A2(n1023), .B1(n1023), .B2(
        uart_phy_rx_phase[13]), .Z(n1024) );
  an02d0 U1670 ( .A1(rs232phy_rs232phyrx_state), .A2(n1024), .Z(N3652) );
  mx02d1 U1671 ( .I0(uart_phy_rx_phase[15]), .I1(n1026), .S(n1025), .Z(n1027)
         );
  an02d0 U1672 ( .A1(n1200), .A2(n1027), .Z(N3654) );
  ah01d1 U1673 ( .A(n1028), .B(uart_phy_tx_phase[12]), .CO(n1030), .S(n1029)
         );
  an02d0 U1674 ( .A1(n2868), .A2(n1029), .Z(N3584) );
  nr03d0 U1675 ( .A1(uart_phy_tx_phase[14]), .A2(uart_phy_tx_phase[13]), .A3(
        n1030), .ZN(n1467) );
  inv0d0 U1676 ( .I(uart_phy_tx_phase[15]), .ZN(n1468) );
  nd02d0 U1677 ( .A1(n1467), .A2(n1468), .ZN(n1128) );
  an02d0 U1678 ( .A1(n2868), .A2(n1031), .Z(N3588) );
  ah01d1 U1679 ( .A(n1032), .B(uart_phy_rx_phase[16]), .CO(n1037), .S(n1033)
         );
  an02d0 U1680 ( .A1(n1200), .A2(n1033), .Z(N3655) );
  an02d0 U1681 ( .A1(mgmtsoc_vexriscv_o_resetOut), .A2(n4881), .Z(N5281) );
  an02d0 U1682 ( .A1(mgmtsoc_vexriscv_reset_debug_logic), .A2(n5956), .Z(N5235) );
  an02d0 U1683 ( .A1(mgmtsoc_litespisdrphycore_posedge_reg), .A2(n5301), .Z(
        N5454) );
  inv0d0 U1684 ( .I(uart_phy_rx_phase[18]), .ZN(n1035) );
  nr02d0 U1685 ( .A1(uart_phy_rx_phase[17]), .A2(n1037), .ZN(n1034) );
  mx02d1 U1686 ( .I0(uart_phy_rx_phase[18]), .I1(n1035), .S(n1034), .Z(n1036)
         );
  an02d0 U1687 ( .A1(n1200), .A2(n1036), .Z(N3657) );
  inv0d0 U1688 ( .I(n1037), .ZN(n1038) );
  aoim22d1 U1689 ( .A1(uart_phy_rx_phase[17]), .A2(n1038), .B1(n1038), .B2(
        uart_phy_rx_phase[17]), .Z(n1039) );
  an02d0 U1690 ( .A1(rs232phy_rs232phyrx_state), .A2(n1039), .Z(N3656) );
  buffd1 U1691 ( .I(n1163), .Z(n1271) );
  nr02d0 U1692 ( .A1(dbg_uart_rx_phase[1]), .A2(dbg_uart_rx_phase[0]), .ZN(
        n1052) );
  inv0d0 U1693 ( .I(dbg_uart_rx_phase[2]), .ZN(n1053) );
  nd02d0 U1694 ( .A1(n1052), .A2(n1053), .ZN(n1066) );
  nr02d0 U1695 ( .A1(dbg_uart_rx_phase[7]), .A2(n1041), .ZN(n1055) );
  inv0d0 U1696 ( .I(dbg_uart_rx_phase[8]), .ZN(n1056) );
  nd02d0 U1697 ( .A1(n1055), .A2(n1056), .ZN(n1046) );
  an02d0 U1698 ( .A1(n1271), .A2(n1040), .Z(N5055) );
  buffd1 U1699 ( .I(n1163), .Z(n1278) );
  inv0d0 U1700 ( .I(n1041), .ZN(n1042) );
  aoim22d1 U1701 ( .A1(dbg_uart_rx_phase[7]), .A2(n1042), .B1(n1042), .B2(
        dbg_uart_rx_phase[7]), .Z(n1043) );
  an02d0 U1702 ( .A1(n1278), .A2(n1043), .Z(N5053) );
  ah01d1 U1703 ( .A(n1044), .B(dbg_uart_rx_phase[4]), .CO(n1064), .S(n1045) );
  an02d0 U1704 ( .A1(n1278), .A2(n1045), .Z(N5050) );
  inv0d0 U1705 ( .I(dbg_uart_rx_phase[12]), .ZN(n1048) );
  ah01d1 U1706 ( .A(n1046), .B(dbg_uart_rx_phase[9]), .CO(n1068), .S(n1040) );
  nr02d0 U1707 ( .A1(dbg_uart_rx_phase[11]), .A2(n1061), .ZN(n1047) );
  mx02d1 U1708 ( .I0(dbg_uart_rx_phase[12]), .I1(n1048), .S(n1047), .Z(n1049)
         );
  an02d0 U1709 ( .A1(n1271), .A2(n1049), .Z(N5058) );
  inv0d0 U1710 ( .I(dbg_uart_rx_phase[0]), .ZN(n1058) );
  an02d0 U1711 ( .A1(n1278), .A2(n1058), .Z(N5046) );
  ah01d1 U1712 ( .A(n1050), .B(dbg_uart_rx_phase[6]), .CO(n1041), .S(n1051) );
  an02d0 U1713 ( .A1(n1278), .A2(n1051), .Z(N5052) );
  mx02d1 U1714 ( .I0(dbg_uart_rx_phase[2]), .I1(n1053), .S(n1052), .Z(n1054)
         );
  an02d0 U1715 ( .A1(n1278), .A2(n1054), .Z(N5048) );
  mx02d1 U1716 ( .I0(dbg_uart_rx_phase[8]), .I1(n1056), .S(n1055), .Z(n1057)
         );
  an02d0 U1717 ( .A1(n1271), .A2(n1057), .Z(N5054) );
  aoim22d1 U1718 ( .A1(dbg_uart_rx_phase[1]), .A2(n1058), .B1(n1058), .B2(
        dbg_uart_rx_phase[1]), .Z(n1059) );
  an02d0 U1719 ( .A1(n1278), .A2(n1059), .Z(N5047) );
  nr03d0 U1720 ( .A1(dbg_uart_rx_phase[12]), .A2(dbg_uart_rx_phase[11]), .A3(
        n1061), .ZN(n1070) );
  aoim22d1 U1721 ( .A1(dbg_uart_rx_phase[13]), .A2(n1070), .B1(n1070), .B2(
        dbg_uart_rx_phase[13]), .Z(n1060) );
  an02d0 U1722 ( .A1(n1271), .A2(n1060), .Z(N5059) );
  inv0d0 U1723 ( .I(n1061), .ZN(n1062) );
  aoim22d1 U1724 ( .A1(dbg_uart_rx_phase[11]), .A2(n1062), .B1(n1062), .B2(
        dbg_uart_rx_phase[11]), .Z(n1063) );
  an02d0 U1725 ( .A1(n1271), .A2(n1063), .Z(N5057) );
  ah01d1 U1726 ( .A(n1064), .B(dbg_uart_rx_phase[5]), .CO(n1050), .S(n1065) );
  an02d0 U1727 ( .A1(n1278), .A2(n1065), .Z(N5051) );
  ah01d1 U1728 ( .A(n1066), .B(dbg_uart_rx_phase[3]), .CO(n1044), .S(n1067) );
  an02d0 U1729 ( .A1(n1278), .A2(n1067), .Z(N5049) );
  ah01d1 U1730 ( .A(n1068), .B(dbg_uart_rx_phase[10]), .CO(n1061), .S(n1069)
         );
  an02d0 U1731 ( .A1(n1271), .A2(n1069), .Z(N5056) );
  inv0d0 U1732 ( .I(dbg_uart_rx_phase[15]), .ZN(n1077) );
  nr02d0 U1733 ( .A1(dbg_uart_rx_phase[14]), .A2(n1072), .ZN(n1078) );
  mx02d1 U1734 ( .I0(dbg_uart_rx_phase[15]), .I1(n1077), .S(n1078), .Z(n1071)
         );
  an02d0 U1735 ( .A1(n1271), .A2(n1071), .Z(N5061) );
  inv0d0 U1736 ( .I(n1072), .ZN(n1073) );
  aoim22d1 U1737 ( .A1(dbg_uart_rx_phase[14]), .A2(n1073), .B1(n1073), .B2(
        dbg_uart_rx_phase[14]), .Z(n1074) );
  an02d0 U1738 ( .A1(n1271), .A2(n1074), .Z(N5060) );
  aoim22d1 U1739 ( .A1(uart_phy_rx_phase[19]), .A2(n1075), .B1(n1075), .B2(
        uart_phy_rx_phase[19]), .Z(n1076) );
  an02d0 U1740 ( .A1(rs232phy_rs232phyrx_state), .A2(n1076), .Z(N3658) );
  nd02d0 U1741 ( .A1(n1078), .A2(n1077), .ZN(n1102) );
  an02d0 U1742 ( .A1(n1271), .A2(n1079), .Z(N5062) );
  nr03d0 U1743 ( .A1(dbg_uart_count[2]), .A2(dbg_uart_count[1]), .A3(
        dbg_uart_count[0]), .ZN(n1091) );
  inv0d0 U1744 ( .I(n1091), .ZN(n1080) );
  nr02d0 U1745 ( .A1(n1080), .A2(dbg_uart_count[3]), .ZN(n1100) );
  inv0d0 U1746 ( .I(dbg_uart_count[5]), .ZN(n1081) );
  aoim22d1 U1747 ( .A1(n1083), .A2(n1081), .B1(n1081), .B2(n1083), .Z(n1082)
         );
  an02d0 U1748 ( .A1(n1171), .A2(n1082), .Z(n4073) );
  nr02d0 U1749 ( .A1(n1083), .A2(dbg_uart_count[5]), .ZN(n2496) );
  nd12d0 U1750 ( .A1(dbg_uart_count[6]), .A2(n2496), .ZN(n1098) );
  nr02d0 U1751 ( .A1(n1098), .A2(dbg_uart_count[7]), .ZN(n1088) );
  aoim22d1 U1752 ( .A1(dbg_uart_count[8]), .A2(n1088), .B1(n1088), .B2(
        dbg_uart_count[8]), .Z(n1084) );
  an02d0 U1753 ( .A1(n1171), .A2(n1084), .Z(n4076) );
  inv0d0 U1754 ( .I(dbg_uart_count[2]), .ZN(n1086) );
  nr02d0 U1755 ( .A1(dbg_uart_count[1]), .A2(dbg_uart_count[0]), .ZN(n1085) );
  mx02d1 U1756 ( .I0(dbg_uart_count[2]), .I1(n1086), .S(n1085), .Z(n1087) );
  an02d0 U1757 ( .A1(n1171), .A2(n1087), .Z(n4070) );
  nr02d0 U1758 ( .A1(n2493), .A2(dbg_uart_count[9]), .ZN(n1093) );
  nd12d0 U1759 ( .A1(dbg_uart_count[10]), .A2(n1093), .ZN(n1111) );
  inv0d0 U1760 ( .I(dbg_uart_count[11]), .ZN(n1089) );
  aoim22d1 U1761 ( .A1(n1111), .A2(n1089), .B1(n1089), .B2(n1111), .Z(n1090)
         );
  an02d0 U1762 ( .A1(n1171), .A2(n1090), .Z(n4079) );
  aoim22d1 U1763 ( .A1(dbg_uart_count[3]), .A2(n1091), .B1(n1091), .B2(
        dbg_uart_count[3]), .Z(n1092) );
  an02d0 U1764 ( .A1(n1171), .A2(n1092), .Z(n4071) );
  aoim22d1 U1765 ( .A1(dbg_uart_count[10]), .A2(n1093), .B1(n1093), .B2(
        dbg_uart_count[10]), .Z(n1094) );
  an02d0 U1766 ( .A1(n1171), .A2(n1094), .Z(n4078) );
  inv0d0 U1767 ( .I(dbg_uart_count[0]), .ZN(n1095) );
  aoim22d1 U1768 ( .A1(dbg_uart_count[1]), .A2(n1095), .B1(n1095), .B2(
        dbg_uart_count[1]), .Z(n1096) );
  an02d0 U1769 ( .A1(n1171), .A2(n1096), .Z(n4069) );
  inv0d0 U1770 ( .I(dbg_uart_count[7]), .ZN(n1097) );
  aoim22d1 U1771 ( .A1(n1098), .A2(n1097), .B1(n1097), .B2(n1098), .Z(n1099)
         );
  an02d0 U1772 ( .A1(n1171), .A2(n1099), .Z(n4075) );
  aoim22d1 U1773 ( .A1(dbg_uart_count[4]), .A2(n1100), .B1(n1100), .B2(
        dbg_uart_count[4]), .Z(n1101) );
  an02d0 U1774 ( .A1(n1171), .A2(n1101), .Z(n4072) );
  ah01d1 U1775 ( .A(n1102), .B(dbg_uart_rx_phase[16]), .CO(n1103), .S(n1079)
         );
  inv0d0 U1776 ( .I(n1103), .ZN(n1130) );
  inv0d0 U1777 ( .I(dbg_uart_rx_phase[17]), .ZN(n1131) );
  aoi22d1 U1778 ( .A1(dbg_uart_rx_phase[17]), .A2(n1130), .B1(n1103), .B2(
        n1131), .ZN(n1104) );
  an02d0 U1779 ( .A1(n1271), .A2(n1104), .Z(N5063) );
  mx02d1 U1780 ( .I0(uart_phy_rx_phase[21]), .I1(n1106), .S(n1105), .Z(n1107)
         );
  an02d0 U1781 ( .A1(n1200), .A2(n1107), .Z(N3660) );
  inv0d0 U1782 ( .I(n1108), .ZN(n1109) );
  aoim22d1 U1783 ( .A1(uart_phy_rx_phase[20]), .A2(n1109), .B1(n1109), .B2(
        uart_phy_rx_phase[20]), .Z(n1110) );
  an02d0 U1784 ( .A1(rs232phy_rs232phyrx_state), .A2(n1110), .Z(N3659) );
  nr02d0 U1785 ( .A1(n1111), .A2(dbg_uart_count[11]), .ZN(n1135) );
  aoim22d1 U1786 ( .A1(dbg_uart_count[12]), .A2(n1135), .B1(n1135), .B2(
        dbg_uart_count[12]), .Z(n1112) );
  an02d0 U1787 ( .A1(n1171), .A2(n1112), .Z(n4080) );
  nd02d0 U1788 ( .A1(uartwishbonebridge_rs232phytx_state), .A2(n4881), .ZN(
        n5990) );
  nr02d0 U1789 ( .A1(dbg_uart_tx_phase[1]), .A2(dbg_uart_tx_phase[0]), .ZN(
        n1719) );
  inv0d0 U1790 ( .I(dbg_uart_tx_phase[2]), .ZN(n1720) );
  nd02d0 U1791 ( .A1(n1719), .A2(n1720), .ZN(n1120) );
  ah01d1 U1792 ( .A(n1114), .B(dbg_uart_tx_phase[5]), .CO(n1116), .S(n1113) );
  ah01d1 U1793 ( .A(n1116), .B(dbg_uart_tx_phase[6]), .CO(n1722), .S(n1115) );
  inv0d0 U1794 ( .I(dbg_uart_tx_phase[8]), .ZN(n1726) );
  nd02d0 U1795 ( .A1(n1725), .A2(n1726), .ZN(n1124) );
  nr03d0 U1796 ( .A1(dbg_uart_tx_phase[12]), .A2(dbg_uart_tx_phase[11]), .A3(
        n1730), .ZN(n1734) );
  nd12d0 U1797 ( .A1(dbg_uart_tx_phase[13]), .A2(n1734), .ZN(n1736) );
  nr02d0 U1798 ( .A1(dbg_uart_tx_phase[14]), .A2(n1736), .ZN(n1739) );
  inv0d0 U1799 ( .I(dbg_uart_tx_phase[15]), .ZN(n1740) );
  nd02d0 U1800 ( .A1(n1739), .A2(n1740), .ZN(n1133) );
  ah01d1 U1801 ( .A(n1118), .B(dbg_uart_tx_phase[4]), .CO(n1114), .S(n1119) );
  ah01d1 U1802 ( .A(n1120), .B(dbg_uart_tx_phase[3]), .CO(n1118), .S(n1121) );
  ah01d1 U1803 ( .A(n1122), .B(dbg_uart_tx_phase[10]), .CO(n1730), .S(n1123)
         );
  ah01d1 U1804 ( .A(n1124), .B(dbg_uart_tx_phase[9]), .CO(n1122), .S(n1125) );
  ah01d1 U1805 ( .A(n1126), .B(uart_phy_rx_phase[22]), .CO(n1140), .S(n1127)
         );
  an02d0 U1806 ( .A1(n1200), .A2(n1127), .Z(N3661) );
  ah01d1 U1807 ( .A(n1128), .B(uart_phy_tx_phase[16]), .CO(n1472), .S(n1031)
         );
  nr03d0 U1808 ( .A1(uart_phy_tx_phase[18]), .A2(uart_phy_tx_phase[17]), .A3(
        n1472), .ZN(n1476) );
  nr02d0 U1809 ( .A1(uart_phy_tx_phase[20]), .A2(n1478), .ZN(n1481) );
  inv0d0 U1810 ( .I(uart_phy_tx_phase[21]), .ZN(n1482) );
  nd02d0 U1811 ( .A1(n1481), .A2(n1482), .ZN(n1138) );
  an02d0 U1812 ( .A1(n2868), .A2(n1129), .Z(N3594) );
  nd02d0 U1813 ( .A1(n1131), .A2(n1130), .ZN(n1142) );
  an02d0 U1814 ( .A1(n1163), .A2(n1132), .Z(N5064) );
  inv0d0 U1815 ( .I(dbg_uart_tx_phase[17]), .ZN(n1742) );
  ah01d1 U1816 ( .A(n1133), .B(dbg_uart_tx_phase[16]), .CO(n1743), .S(n1117)
         );
  inv0d0 U1817 ( .I(n1743), .ZN(n1744) );
  nd02d0 U1818 ( .A1(n1742), .A2(n1744), .ZN(n1144) );
  inv0d0 U1819 ( .I(dbg_uart_count[13]), .ZN(n1136) );
  aoim22d1 U1820 ( .A1(n1168), .A2(n1136), .B1(n1136), .B2(n1168), .Z(n1137)
         );
  an02d0 U1821 ( .A1(n1171), .A2(n1137), .Z(n4081) );
  ah01d1 U1822 ( .A(n1138), .B(uart_phy_tx_phase[22]), .CO(n1148), .S(n1129)
         );
  an02d0 U1823 ( .A1(n2868), .A2(n1139), .Z(N3595) );
  ah01d1 U1824 ( .A(n1140), .B(uart_phy_rx_phase[23]), .CO(n1146), .S(n1141)
         );
  an02d0 U1825 ( .A1(n1200), .A2(n1141), .Z(N3662) );
  ah01d1 U1826 ( .A(n1142), .B(dbg_uart_rx_phase[18]), .CO(n1154), .S(n1132)
         );
  an02d0 U1827 ( .A1(n1278), .A2(n1143), .Z(N5065) );
  ah01d1 U1828 ( .A(n1144), .B(dbg_uart_tx_phase[18]), .CO(n1182), .S(n1134)
         );
  ah01d1 U1829 ( .A(n1146), .B(uart_phy_rx_phase[24]), .CO(n1150), .S(n1147)
         );
  an02d0 U1830 ( .A1(n1200), .A2(n1147), .Z(N3663) );
  ah01d1 U1831 ( .A(n1148), .B(uart_phy_tx_phase[23]), .CO(n1152), .S(n1139)
         );
  an02d0 U1832 ( .A1(n2868), .A2(n1149), .Z(N3596) );
  ah01d1 U1833 ( .A(n1150), .B(uart_phy_rx_phase[25]), .CO(n1164), .S(n1151)
         );
  an02d0 U1834 ( .A1(rs232phy_rs232phyrx_state), .A2(n1151), .Z(N3664) );
  ah01d1 U1835 ( .A(n1152), .B(uart_phy_tx_phase[24]), .CO(n1166), .S(n1149)
         );
  an02d0 U1836 ( .A1(n2868), .A2(n1153), .Z(N3597) );
  inv0d0 U1837 ( .I(dbg_uart_rx_phase[21]), .ZN(n1156) );
  ah01d1 U1838 ( .A(n1154), .B(dbg_uart_rx_phase[19]), .CO(n1172), .S(n1143)
         );
  nr02d0 U1839 ( .A1(dbg_uart_rx_phase[20]), .A2(n1172), .ZN(n1155) );
  mx02d1 U1840 ( .I0(dbg_uart_rx_phase[21]), .I1(n1156), .S(n1155), .Z(n1157)
         );
  an02d0 U1841 ( .A1(n1271), .A2(n1157), .Z(N5067) );
  inv0d0 U1842 ( .I(n1172), .ZN(n1158) );
  aoim22d1 U1843 ( .A1(dbg_uart_rx_phase[20]), .A2(n1158), .B1(n1158), .B2(
        dbg_uart_rx_phase[20]), .Z(n1159) );
  an02d0 U1844 ( .A1(n1278), .A2(n1159), .Z(N5066) );
  inv0d0 U1845 ( .I(dbg_uart_rx_phase[22]), .ZN(n1161) );
  nr03d0 U1846 ( .A1(dbg_uart_rx_phase[21]), .A2(dbg_uart_rx_phase[20]), .A3(
        n1172), .ZN(n1160) );
  mx02d1 U1847 ( .I0(dbg_uart_rx_phase[22]), .I1(n1161), .S(n1160), .Z(n1162)
         );
  an02d0 U1848 ( .A1(n1163), .A2(n1162), .Z(N5068) );
  ah01d1 U1849 ( .A(n1164), .B(uart_phy_rx_phase[26]), .CO(n1176), .S(n1165)
         );
  an02d0 U1850 ( .A1(rs232phy_rs232phyrx_state), .A2(n1165), .Z(N3665) );
  ah01d1 U1851 ( .A(n1166), .B(uart_phy_tx_phase[25]), .CO(n1174), .S(n1153)
         );
  an02d0 U1852 ( .A1(n2868), .A2(n1167), .Z(N3598) );
  nr02d0 U1853 ( .A1(n1168), .A2(dbg_uart_count[13]), .ZN(n2491) );
  nd12d0 U1854 ( .A1(dbg_uart_count[14]), .A2(n2491), .ZN(n2479) );
  inv0d0 U1855 ( .I(dbg_uart_count[15]), .ZN(n1169) );
  aoim22d1 U1856 ( .A1(n2479), .A2(n1169), .B1(n1169), .B2(n2479), .Z(n1170)
         );
  an02d0 U1857 ( .A1(n1171), .A2(n1170), .Z(n4083) );
  inv0d0 U1858 ( .I(dbg_uart_rx_phase[23]), .ZN(n1184) );
  nr04d0 U1859 ( .A1(dbg_uart_rx_phase[22]), .A2(dbg_uart_rx_phase[21]), .A3(
        dbg_uart_rx_phase[20]), .A4(n1172), .ZN(n1185) );
  mx02d1 U1860 ( .I0(dbg_uart_rx_phase[23]), .I1(n1184), .S(n1185), .Z(n1173)
         );
  an02d0 U1861 ( .A1(n1278), .A2(n1173), .Z(N5069) );
  ah01d1 U1862 ( .A(n1174), .B(uart_phy_tx_phase[26]), .CO(n1180), .S(n1167)
         );
  an02d0 U1863 ( .A1(n2868), .A2(n1175), .Z(N3599) );
  ah01d1 U1864 ( .A(n1176), .B(uart_phy_rx_phase[27]), .CO(n1178), .S(n1177)
         );
  an02d0 U1865 ( .A1(rs232phy_rs232phyrx_state), .A2(n1177), .Z(N3666) );
  ah01d1 U1866 ( .A(n1178), .B(uart_phy_rx_phase[28]), .CO(n1187), .S(n1179)
         );
  an02d0 U1867 ( .A1(n1200), .A2(n1179), .Z(N3667) );
  ah01d1 U1868 ( .A(n1180), .B(uart_phy_tx_phase[27]), .CO(n1189), .S(n1175)
         );
  an02d0 U1869 ( .A1(n2868), .A2(n1181), .Z(N3600) );
  ah01d1 U1870 ( .A(n1182), .B(dbg_uart_tx_phase[19]), .CO(n1751), .S(n1145)
         );
  nr04d0 U1871 ( .A1(dbg_uart_tx_phase[22]), .A2(dbg_uart_tx_phase[21]), .A3(
        dbg_uart_tx_phase[20]), .A4(n1751), .ZN(n1755) );
  inv0d0 U1872 ( .I(dbg_uart_tx_phase[23]), .ZN(n1756) );
  nd02d0 U1873 ( .A1(n1755), .A2(n1756), .ZN(n1234) );
  nd02d0 U1874 ( .A1(n1185), .A2(n1184), .ZN(n1195) );
  an02d0 U1875 ( .A1(n1271), .A2(n1186), .Z(N5070) );
  ah01d1 U1876 ( .A(n1187), .B(uart_phy_rx_phase[29]), .CO(n1191), .S(n1188)
         );
  an02d0 U1877 ( .A1(rs232phy_rs232phyrx_state), .A2(n1188), .Z(N3668) );
  ah01d1 U1878 ( .A(n1189), .B(uart_phy_tx_phase[28]), .CO(n1193), .S(n1181)
         );
  an02d0 U1879 ( .A1(n2868), .A2(n1190), .Z(N3601) );
  ah01d1 U1880 ( .A(n1191), .B(uart_phy_rx_phase[30]), .CO(n1198), .S(n1192)
         );
  an02d0 U1881 ( .A1(rs232phy_rs232phyrx_state), .A2(n1192), .Z(N3669) );
  ah01d1 U1882 ( .A(n1193), .B(uart_phy_tx_phase[29]), .CO(n1201), .S(n1190)
         );
  an02d0 U1883 ( .A1(rs232phy_rs232phytx_state), .A2(n1194), .Z(N3602) );
  ah01d1 U1884 ( .A(n1195), .B(dbg_uart_rx_phase[24]), .CO(n1196), .S(n1186)
         );
  inv0d0 U1885 ( .I(n1196), .ZN(n1236) );
  inv0d0 U1886 ( .I(dbg_uart_rx_phase[25]), .ZN(n1237) );
  aoi22d1 U1887 ( .A1(dbg_uart_rx_phase[25]), .A2(n1236), .B1(n1196), .B2(
        n1237), .ZN(n1197) );
  an02d0 U1888 ( .A1(n1278), .A2(n1197), .Z(N5071) );
  ah01d1 U1889 ( .A(n1198), .B(uart_phy_rx_phase[31]), .CO(n1199), .S(n684) );
  an03d0 U1890 ( .A1(n1200), .A2(n1199), .A3(n5288), .Z(N5703) );
  ah01d1 U1891 ( .A(n1201), .B(uart_phy_tx_phase[30]), .CO(n1203), .S(n1194)
         );
  inv0d1 U1892 ( .I(n5111), .ZN(n5301) );
  an03d0 U1893 ( .A1(n2868), .A2(n1202), .A3(n5301), .Z(N5702) );
  ah01d1 U1894 ( .A(n1203), .B(uart_phy_tx_phase[31]), .CO(n1202), .S(n1204)
         );
  an02d0 U1895 ( .A1(n2868), .A2(n1204), .Z(N3603) );
  inv0d0 U1896 ( .I(n4678), .ZN(n3087) );
  an02d0 U1897 ( .A1(n1206), .A2(n4678), .Z(N5644) );
  ah01d1 U1898 ( .A(spi_master_clk_divider1[0]), .B(spi_master_clk_divider1[1]), .CO(n1215), .S(n1206) );
  an02d0 U1899 ( .A1(n1207), .A2(n4678), .Z(N5647) );
  ah01d1 U1900 ( .A(n1208), .B(spi_master_clk_divider1[4]), .CO(n1210), .S(
        n1207) );
  an02d0 U1901 ( .A1(n1209), .A2(n4678), .Z(N5649) );
  ah01d1 U1902 ( .A(n1210), .B(spi_master_clk_divider1[5]), .CO(n1213), .S(
        n1211) );
  an02d0 U1903 ( .A1(n1211), .A2(n4678), .Z(N5648) );
  inv0d0 U1904 ( .I(spi_master_clk_divider1[0]), .ZN(n1212) );
  an02d0 U1905 ( .A1(n1212), .A2(n4678), .Z(N5643) );
  ah01d1 U1906 ( .A(n1213), .B(spi_master_clk_divider1[6]), .CO(n1239), .S(
        n1209) );
  an02d0 U1907 ( .A1(n1214), .A2(n4678), .Z(N5651) );
  ah01d1 U1908 ( .A(n1215), .B(spi_master_clk_divider1[2]), .CO(n1217), .S(
        n1216) );
  an02d0 U1909 ( .A1(n1216), .A2(n4678), .Z(N5645) );
  ah01d1 U1910 ( .A(n1217), .B(spi_master_clk_divider1[3]), .CO(n1208), .S(
        n1218) );
  an02d0 U1911 ( .A1(n1218), .A2(n4678), .Z(N5646) );
  ah01d1 U1912 ( .A(n1219), .B(spi_master_clk_divider1[8]), .CO(n1221), .S(
        n1214) );
  an02d0 U1913 ( .A1(n1220), .A2(n4678), .Z(N5653) );
  ah01d1 U1914 ( .A(n1221), .B(spi_master_clk_divider1[9]), .CO(n1223), .S(
        n1222) );
  an02d0 U1915 ( .A1(n1222), .A2(n4678), .Z(N5652) );
  ah01d1 U1916 ( .A(n1223), .B(spi_master_clk_divider1[10]), .CO(n1232), .S(
        n1220) );
  an02d0 U1917 ( .A1(n1224), .A2(n4678), .Z(N5656) );
  ah01d1 U1918 ( .A(n1225), .B(spi_master_clk_divider1[13]), .CO(n1227), .S(
        n1224) );
  an02d0 U1919 ( .A1(n1226), .A2(n4678), .Z(N5657) );
  ah01d1 U1920 ( .A(n1227), .B(spi_master_clk_divider1[14]), .CO(n1228), .S(
        n1226) );
  xr02d1 U1921 ( .A1(n1228), .A2(spi_master_clk_divider1[15]), .Z(n1229) );
  an02d0 U1922 ( .A1(n1229), .A2(n4678), .Z(N5658) );
  ah01d1 U1923 ( .A(n1230), .B(spi_master_clk_divider1[12]), .CO(n1225), .S(
        n1231) );
  an02d0 U1924 ( .A1(n1231), .A2(n4678), .Z(N5655) );
  ah01d1 U1925 ( .A(n1232), .B(spi_master_clk_divider1[11]), .CO(n1230), .S(
        n1233) );
  an02d0 U1926 ( .A1(n1233), .A2(n4678), .Z(N5654) );
  inv0d0 U1927 ( .I(dbg_uart_tx_phase[25]), .ZN(n1758) );
  ah01d1 U1928 ( .A(n1234), .B(dbg_uart_tx_phase[24]), .CO(n1759), .S(n1183)
         );
  inv0d0 U1929 ( .I(n1759), .ZN(n1760) );
  nd02d0 U1930 ( .A1(n1758), .A2(n1760), .ZN(n1241) );
  nd02d0 U1931 ( .A1(n1237), .A2(n1236), .ZN(n1243) );
  an02d0 U1932 ( .A1(n1271), .A2(n1238), .Z(N5072) );
  ah01d1 U1933 ( .A(n1239), .B(spi_master_clk_divider1[7]), .CO(n1219), .S(
        n1240) );
  an02d0 U1934 ( .A1(n1240), .A2(n4678), .Z(N5650) );
  ah01d1 U1935 ( .A(n1241), .B(dbg_uart_tx_phase[26]), .CO(n1245), .S(n1235)
         );
  ah01d1 U1936 ( .A(n1243), .B(dbg_uart_rx_phase[26]), .CO(n1247), .S(n1238)
         );
  an02d0 U1937 ( .A1(n1278), .A2(n1244), .Z(N5073) );
  ah01d1 U1938 ( .A(n1245), .B(dbg_uart_tx_phase[27]), .CO(n1267), .S(n1242)
         );
  ah01d1 U1939 ( .A(n1247), .B(dbg_uart_rx_phase[27]), .CO(n1269), .S(n1244)
         );
  an02d0 U1940 ( .A1(n1271), .A2(n1248), .Z(N5074) );
  inv0d0 U1941 ( .I(mgmtsoc_litespisdrphycore_sr_cnt[1]), .ZN(n5917) );
  oai21d1 U1942 ( .B1(mgmtsoc_litespisdrphycore_sr_cnt[0]), .B2(n5922), .A(
        n1249), .ZN(n5915) );
  nr03d0 U1943 ( .A1(mgmtsoc_litespisdrphycore_sr_cnt[0]), .A2(n5922), .A3(
        n1249), .ZN(n5914) );
  aoi21d1 U1944 ( .B1(n5917), .B2(n5915), .A(n5914), .ZN(n5929) );
  cg01d0 U1945 ( .A(mgmtsoc_litespisdrphycore_sr_cnt[2]), .B(n5929), .CI(n5928), .CO(n1250) );
  nr02d0 U1946 ( .A1(n1251), .A2(n1250), .ZN(n5942) );
  inv0d0 U1947 ( .I(mgmtsoc_litespisdrphycore_sr_cnt[3]), .ZN(n5940) );
  nr02d0 U1948 ( .A1(n5942), .A2(n5940), .ZN(n5939) );
  oaim21d1 U1949 ( .B1(n1251), .B2(n1250), .A(n1605), .ZN(n5945) );
  nr02d0 U1950 ( .A1(n5939), .A2(n5945), .ZN(n1257) );
  inv0d0 U1951 ( .I(mgmtsoc_litespisdrphycore_sr_cnt[4]), .ZN(n1256) );
  nr02d0 U1952 ( .A1(n5922), .A2(n5921), .ZN(n5920) );
  cg01d0 U1953 ( .A(n5949), .B(n5938), .CI(n5937), .CO(n1254) );
  inv0d0 U1954 ( .I(n1252), .ZN(n1253) );
  nd02d0 U1955 ( .A1(n1253), .A2(n1254), .ZN(n1261) );
  inv0d0 U1956 ( .I(n5941), .ZN(n5951) );
  oan211d1 U1957 ( .C1(n1254), .C2(n1253), .B(n1261), .A(n5951), .ZN(n1255) );
  aoim31d1 U1958 ( .B1(n5941), .B2(n1257), .B3(n1256), .A(n1255), .ZN(n1258)
         );
  nd02d0 U1959 ( .A1(n1257), .A2(n1256), .ZN(n1264) );
  nd02d0 U1960 ( .A1(n1258), .A2(n1264), .ZN(n3123) );
  nr02d0 U1961 ( .A1(mgmtsoc_litespisdrphycore_sr_cnt[5]), .A2(n1264), .ZN(
        n1263) );
  inv0d0 U1962 ( .I(n1263), .ZN(n1259) );
  aoi31d1 U1963 ( .B1(mgmtsoc_litespisdrphycore_sr_cnt[6]), .B2(n5951), .B3(
        n1259), .A(n5950), .ZN(n1260) );
  or02d0 U1964 ( .A1(mgmtsoc_litespisdrphycore_sr_cnt[6]), .A2(n1259), .Z(
        n5953) );
  nd02d0 U1965 ( .A1(n1260), .A2(n5953), .ZN(n3121) );
  aoi31d1 U1966 ( .B1(n5941), .B2(n1262), .B3(n1261), .A(n5950), .ZN(n1266) );
  aoi31d1 U1967 ( .B1(mgmtsoc_litespisdrphycore_sr_cnt[5]), .B2(n5951), .B3(
        n1264), .A(n1263), .ZN(n1265) );
  nd02d0 U1968 ( .A1(n1266), .A2(n1265), .ZN(n3122) );
  ah01d1 U1969 ( .A(n1267), .B(dbg_uart_tx_phase[28]), .CO(n1272), .S(n1246)
         );
  ah01d1 U1970 ( .A(n1269), .B(dbg_uart_rx_phase[28]), .CO(n1274), .S(n1248)
         );
  an02d0 U1971 ( .A1(n1271), .A2(n1270), .Z(N5075) );
  ah01d1 U1972 ( .A(n1272), .B(dbg_uart_tx_phase[29]), .CO(n1279), .S(n1268)
         );
  ah01d1 U1973 ( .A(n1274), .B(dbg_uart_rx_phase[29]), .CO(n1276), .S(n1270)
         );
  an02d0 U1974 ( .A1(n1278), .A2(n1275), .Z(N5076) );
  ah01d1 U1975 ( .A(n1276), .B(dbg_uart_rx_phase[30]), .CO(n1715), .S(n1275)
         );
  an02d0 U1976 ( .A1(n1278), .A2(n1277), .Z(N5757) );
  ah01d1 U1977 ( .A(n1279), .B(dbg_uart_tx_phase[30]), .CO(n1281), .S(n1273)
         );
  ah01d1 U1978 ( .A(n1281), .B(dbg_uart_tx_phase[31]), .CO(n1280), .S(n1282)
         );
  nd12d0 U1979 ( .A1(count[14]), .A2(n1283), .ZN(n1313) );
  inv0d0 U1980 ( .I(count[15]), .ZN(n1284) );
  aoim22d1 U1981 ( .A1(n1313), .A2(n1284), .B1(n1284), .B2(n1313), .Z(n1285)
         );
  aoim22d1 U1982 ( .A1(count[4]), .A2(n1286), .B1(n1286), .B2(count[4]), .Z(
        n1287) );
  aoim22d1 U1983 ( .A1(count[3]), .A2(n1288), .B1(n1288), .B2(count[3]), .Z(
        n1289) );
  aoim22d1 U1984 ( .A1(count[12]), .A2(n1290), .B1(n1290), .B2(count[12]), .Z(
        n1291) );
  inv0d0 U1985 ( .I(count[11]), .ZN(n1292) );
  aoim22d1 U1986 ( .A1(n1293), .A2(n1292), .B1(n1292), .B2(n1293), .Z(n1294)
         );
  inv0d0 U1987 ( .I(count[5]), .ZN(n1295) );
  aoim22d1 U1988 ( .A1(n1296), .A2(n1295), .B1(n1295), .B2(n1296), .Z(n1297)
         );
  inv0d0 U1989 ( .I(count[0]), .ZN(n1298) );
  aoim22d1 U1990 ( .A1(count[1]), .A2(n1298), .B1(n1298), .B2(count[1]), .Z(
        n1299) );
  inv0d0 U1991 ( .I(count[2]), .ZN(n1301) );
  nr02d0 U1992 ( .A1(count[1]), .A2(count[0]), .ZN(n1300) );
  mx02d1 U1993 ( .I0(count[2]), .I1(n1301), .S(n1300), .Z(n1302) );
  inv0d0 U1994 ( .I(count[13]), .ZN(n1303) );
  aoim22d1 U1995 ( .A1(n1304), .A2(n1303), .B1(n1303), .B2(n1304), .Z(n1305)
         );
  aoim22d1 U1996 ( .A1(count[8]), .A2(n1306), .B1(n1306), .B2(count[8]), .Z(
        n1307) );
  inv0d0 U1997 ( .I(count[7]), .ZN(n1308) );
  aoim22d1 U1998 ( .A1(n1309), .A2(n1308), .B1(n1308), .B2(n1309), .Z(n1310)
         );
  aoim22d1 U1999 ( .A1(count[10]), .A2(n1311), .B1(n1311), .B2(count[10]), .Z(
        n1312) );
  an03d0 U2000 ( .A1(n2466), .A2(n2465), .A3(uart_enabled_o), .Z(N4790) );
  an03d0 U2001 ( .A1(n1982), .A2(n2466), .A3(spi_enabled), .Z(N4516) );
  nr02d0 U2002 ( .A1(n1313), .A2(count[15]), .ZN(n1316) );
  nd12d0 U2003 ( .A1(count[16]), .A2(n1316), .ZN(n1319) );
  nr02d0 U2004 ( .A1(n1319), .A2(count[17]), .ZN(n1321) );
  aoim22d1 U2005 ( .A1(count[18]), .A2(n1321), .B1(n1321), .B2(count[18]), .Z(
        n1315) );
  inv0d0 U2006 ( .I(n1314), .ZN(n1887) );
  or02d0 U2007 ( .A1(n1315), .A2(n1887), .Z(n4535) );
  aoim22d1 U2008 ( .A1(count[16]), .A2(n1316), .B1(n1316), .B2(count[16]), .Z(
        n1317) );
  or02d0 U2009 ( .A1(n1317), .A2(n1887), .Z(n4533) );
  inv0d0 U2010 ( .I(count[17]), .ZN(n1318) );
  aoim22d1 U2011 ( .A1(n1319), .A2(n1318), .B1(n1318), .B2(n1319), .Z(n1320)
         );
  or02d0 U2012 ( .A1(n1320), .A2(n1887), .Z(n4534) );
  inv0d0 U2013 ( .I(n1321), .ZN(n1322) );
  oai21d1 U2014 ( .B1(count[18]), .B2(n1322), .A(count[19]), .ZN(n1323) );
  inv0d0 U2015 ( .I(n1323), .ZN(n1324) );
  or02d0 U2016 ( .A1(n1324), .A2(n1887), .Z(n4536) );
  an04d0 U2017 ( .A1(n2476), .A2(n1325), .A3(n1829), .A4(mprj_wb_iena), .Z(
        N4505) );
  inv0d0 U2018 ( .I(n2470), .ZN(n2475) );
  an04d0 U2019 ( .A1(n2476), .A2(n2475), .A3(n2474), .A4(debug_oeb), .Z(N4152)
         );
  nd02d0 U2020 ( .A1(n2474), .A2(n2465), .ZN(n1966) );
  nr02d0 U2021 ( .A1(n1966), .A2(n2654), .ZN(n1924) );
  an02d0 U2022 ( .A1(n5340), .A2(n1924), .Z(N6270) );
  nr04d0 U2023 ( .A1(n1327), .A2(mprj_adr_o[11]), .A3(mprj_adr_o[12]), .A4(
        n1326), .ZN(n1912) );
  inv0d0 U2024 ( .I(n1912), .ZN(n1952) );
  nr02d0 U2025 ( .A1(n1952), .A2(n2654), .ZN(n1916) );
  an02d0 U2026 ( .A1(n5288), .A2(n1916), .Z(N6280) );
  nr02d0 U2027 ( .A1(n1973), .A2(n2654), .ZN(n1928) );
  an02d0 U2028 ( .A1(n5288), .A2(n1928), .Z(N6265) );
  nd02d0 U2029 ( .A1(n2474), .A2(n1328), .ZN(n1937) );
  nr02d0 U2030 ( .A1(n1937), .A2(n2654), .ZN(n1907) );
  an02d0 U2031 ( .A1(n5301), .A2(n1907), .Z(N6290) );
  aoi22d1 U2032 ( .A1(n5401), .A2(\RAM256/Do0_pre[1][26] ), .B1(n5435), .B2(
        \RAM256/Do0_pre[0][26] ), .ZN(n1334) );
  nr04d0 U2033 ( .A1(interface0_bank_bus_dat_r[26]), .A2(
        interface3_bank_bus_dat_r[26]), .A3(interface6_bank_bus_dat_r[26]), 
        .A4(interface10_bank_bus_dat_r[26]), .ZN(n1331) );
  aoi22d1 U2034 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[26]), .B1(slave_sel_r[5]), .B2(hk_dat_i[26]), .ZN(n1330) );
  aoi22d1 U2035 ( .A1(slave_sel_r[0]), .A2(
        mgmtsoc_vexriscv_debug_bus_dat_r[26]), .B1(slave_sel_r[2]), .B2(
        dff2_bus_dat_r[26]), .ZN(n1329) );
  oai211d1 U2036 ( .C1(n1331), .C2(n5356), .A(n1330), .B(n1329), .ZN(n1332) );
  aoi211d1 U2037 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[2]), .C2(
        n1459), .A(n5335), .B(n1332), .ZN(n1333) );
  nd02d0 U2038 ( .A1(n1334), .A2(n1333), .ZN(mgmtsoc_ibus_ibus_dat_r[26]) );
  aoi22d1 U2039 ( .A1(n5437), .A2(\RAM256/Do0_pre[1][18] ), .B1(n1409), .B2(
        \RAM256/Do0_pre[0][18] ), .ZN(n1340) );
  nr04d0 U2040 ( .A1(interface0_bank_bus_dat_r[18]), .A2(
        interface3_bank_bus_dat_r[18]), .A3(interface6_bank_bus_dat_r[18]), 
        .A4(interface10_bank_bus_dat_r[18]), .ZN(n1337) );
  aoi22d1 U2041 ( .A1(n5395), .A2(mgmtsoc_vexriscv_debug_bus_dat_r[18]), .B1(
        slave_sel_r[5]), .B2(hk_dat_i[18]), .ZN(n1336) );
  aoi22d1 U2042 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[18]), .B1(n5406), .B2(
        dff2_bus_dat_r[18]), .ZN(n1335) );
  oai211d1 U2043 ( .C1(n1337), .C2(n5426), .A(n1336), .B(n1335), .ZN(n1338) );
  aoi211d1 U2044 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[10]), 
        .C2(n1459), .A(n1451), .B(n1338), .ZN(n1339) );
  nd02d0 U2045 ( .A1(n1340), .A2(n1339), .ZN(mgmtsoc_ibus_ibus_dat_r[18]) );
  aoi22d1 U2046 ( .A1(n4998), .A2(csrbank10_load0_w[0]), .B1(n1839), .B2(
        csrbank10_value_w[0]), .ZN(n1344) );
  aoi22d1 U2047 ( .A1(n1838), .A2(csrbank10_update_value0_w), .B1(n1806), .B2(
        mgmtsoc_zero1), .ZN(n1343) );
  inv0d0 U2048 ( .I(n1786), .ZN(n4873) );
  aoi22d1 U2049 ( .A1(n1902), .A2(n1614), .B1(n4873), .B2(mgmtsoc_zero2), .ZN(
        n1342) );
  aoi22d1 U2050 ( .A1(n4952), .A2(csrbank10_en0_w), .B1(n2457), .B2(
        csrbank10_reload0_w[0]), .ZN(n1341) );
  an02d0 U2051 ( .A1(n1794), .A2(n1345), .Z(N4694) );
  or02d0 U2052 ( .A1(interface10_bank_bus_dat_r[15]), .A2(
        interface9_bank_bus_dat_r[15]), .Z(n1346) );
  nr04d0 U2053 ( .A1(interface0_bank_bus_dat_r[15]), .A2(
        interface6_bank_bus_dat_r[15]), .A3(interface3_bank_bus_dat_r[15]), 
        .A4(n1346), .ZN(n1349) );
  aoi22d1 U2054 ( .A1(n5394), .A2(mprj_dat_i[15]), .B1(slave_sel_r[0]), .B2(
        mgmtsoc_vexriscv_debug_bus_dat_r[15]), .ZN(n1348) );
  aoi22d1 U2055 ( .A1(n5429), .A2(hk_dat_i[15]), .B1(slave_sel_r[2]), .B2(
        dff2_bus_dat_r[15]), .ZN(n1347) );
  oai211d1 U2056 ( .C1(n1349), .C2(n5426), .A(n1348), .B(n1347), .ZN(n1350) );
  aoi211d1 U2057 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[23]), 
        .C2(n1459), .A(n1451), .B(n1350), .ZN(n1352) );
  aoi22d1 U2058 ( .A1(n5401), .A2(\RAM256/Do0_pre[1][15] ), .B1(n1409), .B2(
        \RAM256/Do0_pre[0][15] ), .ZN(n1351) );
  nd02d0 U2059 ( .A1(n1352), .A2(n1351), .ZN(mgmtsoc_ibus_ibus_dat_r[15]) );
  aoi22d1 U2060 ( .A1(n5401), .A2(\RAM256/Do0_pre[1][21] ), .B1(n5435), .B2(
        \RAM256/Do0_pre[0][21] ), .ZN(n1358) );
  nr04d0 U2061 ( .A1(interface0_bank_bus_dat_r[21]), .A2(
        interface3_bank_bus_dat_r[21]), .A3(interface6_bank_bus_dat_r[21]), 
        .A4(interface10_bank_bus_dat_r[21]), .ZN(n1355) );
  aoi22d1 U2062 ( .A1(slave_sel_r[0]), .A2(
        mgmtsoc_vexriscv_debug_bus_dat_r[21]), .B1(slave_sel_r[5]), .B2(
        hk_dat_i[21]), .ZN(n1354) );
  aoi22d1 U2063 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[21]), .B1(slave_sel_r[2]), .B2(dff2_bus_dat_r[21]), .ZN(n1353) );
  oai211d1 U2064 ( .C1(n1355), .C2(n5426), .A(n1354), .B(n1353), .ZN(n1356) );
  aoi211d1 U2065 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[13]), 
        .C2(n1459), .A(n1451), .B(n1356), .ZN(n1357) );
  nd02d0 U2066 ( .A1(n1358), .A2(n1357), .ZN(mgmtsoc_ibus_ibus_dat_r[21]) );
  aoi22d1 U2067 ( .A1(n5401), .A2(\RAM256/Do0_pre[1][17] ), .B1(n5435), .B2(
        \RAM256/Do0_pre[0][17] ), .ZN(n1364) );
  nr04d0 U2068 ( .A1(interface0_bank_bus_dat_r[17]), .A2(
        interface3_bank_bus_dat_r[17]), .A3(interface6_bank_bus_dat_r[17]), 
        .A4(interface10_bank_bus_dat_r[17]), .ZN(n1361) );
  aoi22d1 U2069 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[17]), .B1(slave_sel_r[2]), .B2(dff2_bus_dat_r[17]), .ZN(n1360) );
  aoi22d1 U2070 ( .A1(n5395), .A2(mgmtsoc_vexriscv_debug_bus_dat_r[17]), .B1(
        n5429), .B2(hk_dat_i[17]), .ZN(n1359) );
  oai211d1 U2071 ( .C1(n1361), .C2(n5356), .A(n1360), .B(n1359), .ZN(n1362) );
  aoi211d1 U2072 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[9]), .C2(
        n1459), .A(n1451), .B(n1362), .ZN(n1363) );
  nd02d0 U2073 ( .A1(n1364), .A2(n1363), .ZN(mgmtsoc_ibus_ibus_dat_r[17]) );
  aoi22d1 U2074 ( .A1(n5401), .A2(\RAM256/Do0_pre[1][28] ), .B1(n1409), .B2(
        \RAM256/Do0_pre[0][28] ), .ZN(n1370) );
  nr04d0 U2075 ( .A1(interface0_bank_bus_dat_r[28]), .A2(
        interface3_bank_bus_dat_r[28]), .A3(interface6_bank_bus_dat_r[28]), 
        .A4(interface10_bank_bus_dat_r[28]), .ZN(n1367) );
  aoi22d1 U2076 ( .A1(n5394), .A2(mprj_dat_i[28]), .B1(n5395), .B2(
        mgmtsoc_vexriscv_debug_bus_dat_r[28]), .ZN(n1366) );
  aoi22d1 U2077 ( .A1(n5429), .A2(hk_dat_i[28]), .B1(n5406), .B2(
        dff2_bus_dat_r[28]), .ZN(n1365) );
  oai211d1 U2078 ( .C1(n1367), .C2(n5356), .A(n1366), .B(n1365), .ZN(n1368) );
  aoi211d1 U2079 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[4]), .C2(
        n1459), .A(n5335), .B(n1368), .ZN(n1369) );
  nd02d0 U2080 ( .A1(n1370), .A2(n1369), .ZN(mgmtsoc_ibus_ibus_dat_r[28]) );
  aoi22d1 U2081 ( .A1(n5401), .A2(\RAM256/Do0_pre[1][31] ), .B1(n1409), .B2(
        \RAM256/Do0_pre[0][31] ), .ZN(n1376) );
  nr04d0 U2082 ( .A1(interface0_bank_bus_dat_r[31]), .A2(
        interface3_bank_bus_dat_r[31]), .A3(interface6_bank_bus_dat_r[31]), 
        .A4(interface10_bank_bus_dat_r[31]), .ZN(n1373) );
  aoi22d1 U2083 ( .A1(n5394), .A2(mprj_dat_i[31]), .B1(slave_sel_r[5]), .B2(
        hk_dat_i[31]), .ZN(n1372) );
  aoi22d1 U2084 ( .A1(slave_sel_r[0]), .A2(
        mgmtsoc_vexriscv_debug_bus_dat_r[31]), .B1(n5406), .B2(
        dff2_bus_dat_r[31]), .ZN(n1371) );
  oai211d1 U2085 ( .C1(n1373), .C2(n5356), .A(n1372), .B(n1371), .ZN(n1374) );
  aoi211d1 U2086 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[7]), .C2(
        n1459), .A(n1451), .B(n1374), .ZN(n1375) );
  nd02d0 U2087 ( .A1(n1376), .A2(n1375), .ZN(mgmtsoc_ibus_ibus_dat_r[31]) );
  aoi22d1 U2088 ( .A1(n5401), .A2(\RAM256/Do0_pre[1][29] ), .B1(n1409), .B2(
        \RAM256/Do0_pre[0][29] ), .ZN(n1382) );
  aoi22d1 U2089 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[29]), .B1(slave_sel_r[2]), .B2(dff2_bus_dat_r[29]), .ZN(n1378) );
  aoi22d1 U2090 ( .A1(slave_sel_r[0]), .A2(
        mgmtsoc_vexriscv_debug_bus_dat_r[29]), .B1(n5429), .B2(hk_dat_i[29]), 
        .ZN(n1377) );
  oai211d1 U2091 ( .C1(n1379), .C2(n5356), .A(n1378), .B(n1377), .ZN(n1380) );
  aoi211d1 U2092 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[5]), .C2(
        n1459), .A(n5335), .B(n1380), .ZN(n1381) );
  nd02d0 U2093 ( .A1(n1382), .A2(n1381), .ZN(mgmtsoc_ibus_ibus_dat_r[29]) );
  or04d0 U2094 ( .A1(interface9_bank_bus_dat_r[5]), .A2(
        interface10_bank_bus_dat_r[5]), .A3(interface0_bank_bus_dat_r[5]), 
        .A4(interface11_bank_bus_dat_r[5]), .Z(n1383) );
  nr04d0 U2095 ( .A1(interface3_bank_bus_dat_r[5]), .A2(
        interface6_bank_bus_dat_r[5]), .A3(interface4_bank_bus_dat_r[5]), .A4(
        n1383), .ZN(n1386) );
  aoi22d1 U2096 ( .A1(n5394), .A2(mprj_dat_i[5]), .B1(slave_sel_r[0]), .B2(
        mgmtsoc_vexriscv_debug_bus_dat_r[5]), .ZN(n1385) );
  aoi22d1 U2097 ( .A1(n5429), .A2(hk_dat_i[5]), .B1(n5406), .B2(
        dff2_bus_dat_r[5]), .ZN(n1384) );
  oai211d1 U2098 ( .C1(n1386), .C2(n5426), .A(n1385), .B(n1384), .ZN(n1387) );
  aoi211d1 U2099 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[29]), 
        .C2(n1459), .A(n5335), .B(n1387), .ZN(n1389) );
  aoi22d1 U2100 ( .A1(n5437), .A2(\RAM256/Do0_pre[1][5] ), .B1(n5435), .B2(
        \RAM256/Do0_pre[0][5] ), .ZN(n1388) );
  or02d0 U2101 ( .A1(interface10_bank_bus_dat_r[16]), .A2(
        interface9_bank_bus_dat_r[16]), .Z(n1390) );
  nr04d0 U2102 ( .A1(interface0_bank_bus_dat_r[16]), .A2(
        interface6_bank_bus_dat_r[16]), .A3(interface3_bank_bus_dat_r[16]), 
        .A4(n1390), .ZN(n1393) );
  aoi22d1 U2103 ( .A1(n5394), .A2(mprj_dat_i[16]), .B1(slave_sel_r[2]), .B2(
        dff2_bus_dat_r[16]), .ZN(n1392) );
  aoi22d1 U2104 ( .A1(n5395), .A2(mgmtsoc_vexriscv_debug_bus_dat_r[16]), .B1(
        slave_sel_r[5]), .B2(hk_dat_i[16]), .ZN(n1391) );
  oai211d1 U2105 ( .C1(n1393), .C2(n5356), .A(n1392), .B(n1391), .ZN(n1394) );
  aoi211d1 U2106 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[8]), .C2(
        n1459), .A(n1451), .B(n1394), .ZN(n1396) );
  aoi22d1 U2107 ( .A1(n5437), .A2(\RAM256/Do0_pre[1][16] ), .B1(n1409), .B2(
        \RAM256/Do0_pre[0][16] ), .ZN(n1395) );
  nd02d0 U2108 ( .A1(n1396), .A2(n1395), .ZN(mgmtsoc_ibus_ibus_dat_r[16]) );
  aoi22d1 U2109 ( .A1(n5437), .A2(\RAM256/Do0_pre[1][22] ), .B1(n1409), .B2(
        \RAM256/Do0_pre[0][22] ), .ZN(n1402) );
  nr04d0 U2110 ( .A1(interface0_bank_bus_dat_r[22]), .A2(
        interface3_bank_bus_dat_r[22]), .A3(interface6_bank_bus_dat_r[22]), 
        .A4(interface10_bank_bus_dat_r[22]), .ZN(n1399) );
  aoi22d1 U2111 ( .A1(n5394), .A2(mprj_dat_i[22]), .B1(slave_sel_r[2]), .B2(
        dff2_bus_dat_r[22]), .ZN(n1398) );
  aoi22d1 U2112 ( .A1(slave_sel_r[0]), .A2(
        mgmtsoc_vexriscv_debug_bus_dat_r[22]), .B1(n5429), .B2(hk_dat_i[22]), 
        .ZN(n1397) );
  oai211d1 U2113 ( .C1(n1399), .C2(n5356), .A(n1398), .B(n1397), .ZN(n1400) );
  aoi211d1 U2114 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[14]), 
        .C2(n1459), .A(n5335), .B(n1400), .ZN(n1401) );
  nd02d0 U2115 ( .A1(n1402), .A2(n1401), .ZN(mgmtsoc_ibus_ibus_dat_r[22]) );
  aoi22d1 U2116 ( .A1(n5401), .A2(\RAM256/Do0_pre[1][27] ), .B1(n1409), .B2(
        \RAM256/Do0_pre[0][27] ), .ZN(n1408) );
  nr04d0 U2117 ( .A1(interface0_bank_bus_dat_r[27]), .A2(
        interface3_bank_bus_dat_r[27]), .A3(interface6_bank_bus_dat_r[27]), 
        .A4(interface10_bank_bus_dat_r[27]), .ZN(n1405) );
  aoi22d1 U2118 ( .A1(slave_sel_r[0]), .A2(
        mgmtsoc_vexriscv_debug_bus_dat_r[27]), .B1(n5406), .B2(
        dff2_bus_dat_r[27]), .ZN(n1404) );
  aoi22d1 U2119 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[27]), .B1(slave_sel_r[5]), .B2(hk_dat_i[27]), .ZN(n1403) );
  oai211d1 U2120 ( .C1(n1405), .C2(n5356), .A(n1404), .B(n1403), .ZN(n1406) );
  aoi211d1 U2121 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[3]), .C2(
        n1459), .A(n5335), .B(n1406), .ZN(n1407) );
  nd02d0 U2122 ( .A1(n1408), .A2(n1407), .ZN(mgmtsoc_ibus_ibus_dat_r[27]) );
  aoi22d1 U2123 ( .A1(n5437), .A2(\RAM256/Do0_pre[1][20] ), .B1(n1409), .B2(
        \RAM256/Do0_pre[0][20] ), .ZN(n1415) );
  nr04d0 U2124 ( .A1(interface0_bank_bus_dat_r[20]), .A2(
        interface3_bank_bus_dat_r[20]), .A3(interface6_bank_bus_dat_r[20]), 
        .A4(interface10_bank_bus_dat_r[20]), .ZN(n1412) );
  aoi22d1 U2125 ( .A1(slave_sel_r[5]), .A2(hk_dat_i[20]), .B1(slave_sel_r[2]), 
        .B2(dff2_bus_dat_r[20]), .ZN(n1411) );
  aoi22d1 U2126 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[20]), .B1(slave_sel_r[0]), .B2(mgmtsoc_vexriscv_debug_bus_dat_r[20]), .ZN(n1410) );
  oai211d1 U2127 ( .C1(n1412), .C2(n5356), .A(n1411), .B(n1410), .ZN(n1413) );
  aoi211d1 U2128 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[12]), 
        .C2(n1459), .A(n1451), .B(n1413), .ZN(n1414) );
  nd02d0 U2129 ( .A1(n1415), .A2(n1414), .ZN(mgmtsoc_ibus_ibus_dat_r[20]) );
  aoi22d1 U2130 ( .A1(n5401), .A2(\RAM256/Do0_pre[1][30] ), .B1(n5435), .B2(
        \RAM256/Do0_pre[0][30] ), .ZN(n1421) );
  nr04d0 U2131 ( .A1(interface0_bank_bus_dat_r[30]), .A2(
        interface3_bank_bus_dat_r[30]), .A3(interface6_bank_bus_dat_r[30]), 
        .A4(interface10_bank_bus_dat_r[30]), .ZN(n1418) );
  aoi22d1 U2132 ( .A1(n5429), .A2(hk_dat_i[30]), .B1(slave_sel_r[2]), .B2(
        dff2_bus_dat_r[30]), .ZN(n1417) );
  aoi22d1 U2133 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[30]), .B1(n5395), .B2(
        mgmtsoc_vexriscv_debug_bus_dat_r[30]), .ZN(n1416) );
  oai211d1 U2134 ( .C1(n1418), .C2(n5356), .A(n1417), .B(n1416), .ZN(n1419) );
  aoi211d1 U2135 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[6]), .C2(
        n1459), .A(n5335), .B(n1419), .ZN(n1420) );
  nd02d0 U2136 ( .A1(n1421), .A2(n1420), .ZN(mgmtsoc_ibus_ibus_dat_r[30]) );
  aoi22d1 U2137 ( .A1(n5401), .A2(\RAM256/Do0_pre[1][25] ), .B1(n5435), .B2(
        \RAM256/Do0_pre[0][25] ), .ZN(n1427) );
  nr04d0 U2138 ( .A1(interface0_bank_bus_dat_r[25]), .A2(
        interface3_bank_bus_dat_r[25]), .A3(interface6_bank_bus_dat_r[25]), 
        .A4(interface10_bank_bus_dat_r[25]), .ZN(n1424) );
  aoi22d1 U2139 ( .A1(n5394), .A2(mprj_dat_i[25]), .B1(n5395), .B2(
        mgmtsoc_vexriscv_debug_bus_dat_r[25]), .ZN(n1423) );
  aoi22d1 U2140 ( .A1(slave_sel_r[5]), .A2(hk_dat_i[25]), .B1(slave_sel_r[2]), 
        .B2(dff2_bus_dat_r[25]), .ZN(n1422) );
  oai211d1 U2141 ( .C1(n1424), .C2(n5426), .A(n1423), .B(n1422), .ZN(n1425) );
  aoi211d1 U2142 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[1]), .C2(
        n1459), .A(n5335), .B(n1425), .ZN(n1426) );
  nd02d0 U2143 ( .A1(n1427), .A2(n1426), .ZN(mgmtsoc_ibus_ibus_dat_r[25]) );
  aoi22d1 U2144 ( .A1(n5401), .A2(\RAM256/Do0_pre[1][24] ), .B1(n5435), .B2(
        \RAM256/Do0_pre[0][24] ), .ZN(n1433) );
  aoi22d1 U2145 ( .A1(n5429), .A2(hk_dat_i[24]), .B1(slave_sel_r[2]), .B2(
        dff2_bus_dat_r[24]), .ZN(n1429) );
  aoi22d1 U2146 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[24]), .B1(slave_sel_r[0]), .B2(mgmtsoc_vexriscv_debug_bus_dat_r[24]), .ZN(n1428) );
  oai211d1 U2147 ( .C1(n1430), .C2(n5426), .A(n1429), .B(n1428), .ZN(n1431) );
  aoi211d1 U2148 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[0]), .C2(
        n1459), .A(n5335), .B(n1431), .ZN(n1432) );
  nd02d0 U2149 ( .A1(n1433), .A2(n1432), .ZN(mgmtsoc_ibus_ibus_dat_r[24]) );
  aoi22d1 U2150 ( .A1(n5401), .A2(\RAM256/Do0_pre[1][23] ), .B1(n1409), .B2(
        \RAM256/Do0_pre[0][23] ), .ZN(n1439) );
  nr04d0 U2151 ( .A1(interface0_bank_bus_dat_r[23]), .A2(
        interface3_bank_bus_dat_r[23]), .A3(interface6_bank_bus_dat_r[23]), 
        .A4(interface10_bank_bus_dat_r[23]), .ZN(n1436) );
  aoi22d1 U2152 ( .A1(n5395), .A2(mgmtsoc_vexriscv_debug_bus_dat_r[23]), .B1(
        slave_sel_r[5]), .B2(hk_dat_i[23]), .ZN(n1435) );
  aoi22d1 U2153 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[23]), .B1(n5406), .B2(
        dff2_bus_dat_r[23]), .ZN(n1434) );
  oai211d1 U2154 ( .C1(n1436), .C2(n5426), .A(n1435), .B(n1434), .ZN(n1437) );
  aoi211d1 U2155 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[15]), 
        .C2(n1459), .A(n5335), .B(n1437), .ZN(n1438) );
  nd02d0 U2156 ( .A1(n1439), .A2(n1438), .ZN(mgmtsoc_ibus_ibus_dat_r[23]) );
  aoi22d1 U2157 ( .A1(n5401), .A2(\RAM256/Do0_pre[1][19] ), .B1(n1409), .B2(
        \RAM256/Do0_pre[0][19] ), .ZN(n1445) );
  aoi22d1 U2158 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[19]), .B1(slave_sel_r[2]), .B2(dff2_bus_dat_r[19]), .ZN(n1441) );
  aoi22d1 U2159 ( .A1(n5395), .A2(mgmtsoc_vexriscv_debug_bus_dat_r[19]), .B1(
        slave_sel_r[5]), .B2(hk_dat_i[19]), .ZN(n1440) );
  oai211d1 U2160 ( .C1(n1442), .C2(n5356), .A(n1441), .B(n1440), .ZN(n1443) );
  aoi211d1 U2161 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[11]), 
        .C2(n1459), .A(n1451), .B(n1443), .ZN(n1444) );
  nd02d0 U2162 ( .A1(n1445), .A2(n1444), .ZN(mgmtsoc_ibus_ibus_dat_r[19]) );
  or02d0 U2163 ( .A1(interface10_bank_bus_dat_r[12]), .A2(
        interface9_bank_bus_dat_r[12]), .Z(n1446) );
  nr04d0 U2164 ( .A1(interface0_bank_bus_dat_r[12]), .A2(
        interface6_bank_bus_dat_r[12]), .A3(interface3_bank_bus_dat_r[12]), 
        .A4(n1446), .ZN(n1449) );
  aoi22d1 U2165 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[12]), .B1(n5395), .B2(
        mgmtsoc_vexriscv_debug_bus_dat_r[12]), .ZN(n1448) );
  aoi22d1 U2166 ( .A1(n5429), .A2(hk_dat_i[12]), .B1(slave_sel_r[2]), .B2(
        dff2_bus_dat_r[12]), .ZN(n1447) );
  oai211d1 U2167 ( .C1(n1449), .C2(n5426), .A(n1448), .B(n1447), .ZN(n1450) );
  aoi211d1 U2168 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[20]), 
        .C2(n1459), .A(n1451), .B(n1450), .ZN(n1453) );
  aoi22d1 U2169 ( .A1(n5437), .A2(\RAM256/Do0_pre[1][12] ), .B1(n5435), .B2(
        \RAM256/Do0_pre[0][12] ), .ZN(n1452) );
  nd02d0 U2170 ( .A1(n1453), .A2(n1452), .ZN(mgmtsoc_ibus_ibus_dat_r[12]) );
  or04d0 U2171 ( .A1(interface9_bank_bus_dat_r[4]), .A2(
        interface10_bank_bus_dat_r[4]), .A3(interface0_bank_bus_dat_r[4]), 
        .A4(interface11_bank_bus_dat_r[4]), .Z(n1454) );
  nr04d0 U2172 ( .A1(interface3_bank_bus_dat_r[4]), .A2(
        interface6_bank_bus_dat_r[4]), .A3(interface4_bank_bus_dat_r[4]), .A4(
        n1454), .ZN(n1457) );
  aoi22d1 U2173 ( .A1(n5394), .A2(mprj_dat_i[4]), .B1(n5395), .B2(
        mgmtsoc_vexriscv_debug_bus_dat_r[4]), .ZN(n1456) );
  aoi22d1 U2174 ( .A1(n5429), .A2(hk_dat_i[4]), .B1(n5406), .B2(
        dff2_bus_dat_r[4]), .ZN(n1455) );
  oai211d1 U2175 ( .C1(n1457), .C2(n5426), .A(n1456), .B(n1455), .ZN(n1458) );
  aoi211d1 U2176 ( .C1(mgmtsoc_litespisdrphycore_source_payload_data[28]), 
        .C2(n1459), .A(n5335), .B(n1458), .ZN(n1461) );
  aoi22d1 U2177 ( .A1(n5437), .A2(\RAM256/Do0_pre[1][4] ), .B1(n5435), .B2(
        \RAM256/Do0_pre[0][4] ), .ZN(n1460) );
  nd02d0 U2178 ( .A1(n1461), .A2(n1460), .ZN(mgmtsoc_ibus_ibus_dat_r[4]) );
  aor22d1 U2180 ( .A1(csrbank11_ev_enable0_w[0]), .A2(uart_pending_status[0]), 
        .B1(csrbank11_ev_enable0_w[1]), .B2(uart_pending_status[1]), .Z(
        mgmtsoc_interrupt[1]) );
  inv0d0 U2181 ( .I(uart_phy_tx_phase[5]), .ZN(n1462) );
  nd12d0 U2182 ( .A1(n1462), .A2(rs232phy_rs232phytx_state), .ZN(N3577) );
  aoi22d1 U2183 ( .A1(uart_phy_tx_phase[9]), .A2(n1465), .B1(n1464), .B2(n1463), .ZN(n1466) );
  nd12d0 U2184 ( .A1(n1466), .A2(rs232phy_rs232phytx_state), .ZN(N3581) );
  mx02d1 U2185 ( .I0(uart_phy_tx_phase[15]), .I1(n1468), .S(n1467), .Z(n1469)
         );
  nd12d0 U2186 ( .A1(n1469), .A2(rs232phy_rs232phytx_state), .ZN(N3587) );
  inv0d0 U2187 ( .I(n1472), .ZN(n1470) );
  aoim22d1 U2188 ( .A1(uart_phy_tx_phase[17]), .A2(n1470), .B1(n1470), .B2(
        uart_phy_tx_phase[17]), .Z(n1471) );
  nd12d0 U2189 ( .A1(n1471), .A2(rs232phy_rs232phytx_state), .ZN(N3589) );
  inv0d0 U2190 ( .I(uart_phy_tx_phase[18]), .ZN(n1474) );
  nr02d0 U2191 ( .A1(uart_phy_tx_phase[17]), .A2(n1472), .ZN(n1473) );
  mx02d1 U2192 ( .I0(uart_phy_tx_phase[18]), .I1(n1474), .S(n1473), .Z(n1475)
         );
  nd12d0 U2193 ( .A1(n1475), .A2(rs232phy_rs232phytx_state), .ZN(N3590) );
  aoim22d1 U2194 ( .A1(uart_phy_tx_phase[19]), .A2(n1476), .B1(n1476), .B2(
        uart_phy_tx_phase[19]), .Z(n1477) );
  nd12d0 U2195 ( .A1(n1477), .A2(rs232phy_rs232phytx_state), .ZN(N3591) );
  inv0d0 U2196 ( .I(n1478), .ZN(n1479) );
  aoim22d1 U2197 ( .A1(uart_phy_tx_phase[20]), .A2(n1479), .B1(n1479), .B2(
        uart_phy_tx_phase[20]), .Z(n1480) );
  nd12d0 U2198 ( .A1(n1480), .A2(rs232phy_rs232phytx_state), .ZN(N3592) );
  mx02d1 U2199 ( .I0(uart_phy_tx_phase[21]), .I1(n1482), .S(n1481), .Z(n1483)
         );
  nd12d0 U2200 ( .A1(n1483), .A2(rs232phy_rs232phytx_state), .ZN(N3593) );
  inv0d0 U2201 ( .I(dbg_uart_length[5]), .ZN(n1484) );
  nr03d0 U2202 ( .A1(dbg_uart_length[2]), .A2(dbg_uart_length[1]), .A3(
        dbg_uart_length[0]), .ZN(n1488) );
  inv0d0 U2203 ( .I(dbg_uart_length[3]), .ZN(n1486) );
  nd02d0 U2204 ( .A1(n1488), .A2(n1486), .ZN(n1493) );
  inv0d0 U2205 ( .I(dbg_uart_length[4]), .ZN(n1494) );
  nd12d0 U2206 ( .A1(n1493), .A2(n1494), .ZN(n1502) );
  mx02d1 U2207 ( .I0(dbg_uart_length[5]), .I1(n1484), .S(n1502), .Z(n1501) );
  inv0d0 U2208 ( .I(dbg_uart_length[2]), .ZN(n1485) );
  mx02d1 U2209 ( .I0(n1485), .I1(dbg_uart_length[2]), .S(
        dbg_uart_words_count[2]), .Z(n1491) );
  nr02d0 U2210 ( .A1(dbg_uart_length[1]), .A2(dbg_uart_length[0]), .ZN(n1490)
         );
  mx02d1 U2211 ( .I0(n1486), .I1(dbg_uart_length[3]), .S(
        dbg_uart_words_count[3]), .Z(n1489) );
  oai22d1 U2212 ( .A1(n1488), .A2(n1489), .B1(n1490), .B2(n1491), .ZN(n1487)
         );
  aoi221d1 U2213 ( .B1(n1491), .B2(n1490), .C1(n1489), .C2(n1488), .A(n1487), 
        .ZN(n1500) );
  inv0d0 U2214 ( .I(dbg_uart_length[1]), .ZN(n1492) );
  mx02d1 U2215 ( .I0(n1492), .I1(dbg_uart_length[1]), .S(
        dbg_uart_words_count[1]), .Z(n1497) );
  xr03d1 U2216 ( .A1(n1494), .A2(n1493), .A3(dbg_uart_words_count[4]), .Z(
        n1495) );
  oan211d1 U2217 ( .C1(dbg_uart_length[0]), .C2(n1497), .B(
        dbg_uart_words_count[0]), .A(n1495), .ZN(n1496) );
  aon211d1 U2218 ( .C1(dbg_uart_length[0]), .C2(n1497), .B(
        dbg_uart_words_count[0]), .A(n1496), .ZN(n1498) );
  aoi21d1 U2219 ( .B1(n1501), .B2(dbg_uart_words_count[5]), .A(n1498), .ZN(
        n1499) );
  oai211d1 U2220 ( .C1(n1501), .C2(dbg_uart_words_count[5]), .A(n1500), .B(
        n1499), .ZN(n1512) );
  nr02d0 U2221 ( .A1(dbg_uart_length[5]), .A2(n1502), .ZN(n1504) );
  inv0d0 U2222 ( .I(dbg_uart_length[6]), .ZN(n1503) );
  nd02d0 U2223 ( .A1(n1504), .A2(n1503), .ZN(n1510) );
  nr02d0 U2224 ( .A1(n1504), .A2(n1503), .ZN(n1505) );
  inv0d0 U2225 ( .I(n1505), .ZN(n1509) );
  xr02d1 U2226 ( .A1(dbg_uart_length[7]), .A2(dbg_uart_words_count[7]), .Z(
        n1506) );
  nr02d0 U2227 ( .A1(n1505), .A2(n1506), .ZN(n1507) );
  aoi22d1 U2228 ( .A1(dbg_uart_words_count[6]), .A2(n1507), .B1(n1506), .B2(
        n1510), .ZN(n1508) );
  aon211d1 U2229 ( .C1(n1510), .C2(n1509), .B(dbg_uart_words_count[6]), .A(
        n1508), .ZN(n1511) );
  nr02d0 U2230 ( .A1(n1512), .A2(n1511), .ZN(n1525) );
  inv0d0 U2231 ( .I(n1525), .ZN(n1536) );
  nd03d0 U2232 ( .A1(uartwishbonebridge_state[1]), .A2(
        uartwishbonebridge_state[2]), .A3(n5488), .ZN(n5300) );
  nd02d0 U2233 ( .A1(dbg_uart_bytes_count[0]), .A2(dbg_uart_bytes_count[1]), 
        .ZN(n5986) );
  nd02d0 U2234 ( .A1(dbg_uart_tx_tick), .A2(dbg_uart_tx_count[0]), .ZN(n5979)
         );
  inv0d0 U2235 ( .I(dbg_uart_tx_count[3]), .ZN(n5984) );
  nr04d0 U2236 ( .A1(dbg_uart_tx_count[1]), .A2(dbg_uart_tx_count[2]), .A3(
        n5979), .A4(n5984), .ZN(n5985) );
  nd02d0 U2237 ( .A1(uartwishbonebridge_rs232phytx_state), .A2(n5985), .ZN(
        n1535) );
  inv0d0 U2238 ( .I(n1522), .ZN(n5299) );
  oai22d1 U2239 ( .A1(n1513), .A2(n1532), .B1(n5300), .B2(n5299), .ZN(n5491)
         );
  inv0d0 U2240 ( .I(n1524), .ZN(n1516) );
  nr02d0 U2241 ( .A1(uartwishbonebridge_state[2]), .A2(n5296), .ZN(n5489) );
  nr02d0 U2242 ( .A1(n5986), .A2(n5342), .ZN(n1538) );
  inv0d0 U2243 ( .I(n5341), .ZN(n1527) );
  nr04d0 U2244 ( .A1(n1529), .A2(n1538), .A3(n1527), .A4(n5488), .ZN(n1517) );
  nd02d0 U2245 ( .A1(n2482), .A2(n1516), .ZN(n5954) );
  inv0d0 U2246 ( .I(n5954), .ZN(n5957) );
  aoi211d1 U2247 ( .C1(n1536), .C2(n5491), .A(n1517), .B(n5957), .ZN(n1521) );
  nd02d0 U2248 ( .A1(n1538), .A2(n5488), .ZN(n2506) );
  nr02d0 U2249 ( .A1(n2504), .A2(n2506), .ZN(n1520) );
  inv0d0 U2250 ( .I(dbg_uart_cmd[7]), .ZN(n5967) );
  inv0d0 U2251 ( .I(dbg_uart_cmd[6]), .ZN(n5964) );
  nd02d0 U2252 ( .A1(n5967), .A2(n5964), .ZN(n1518) );
  nr04d0 U2253 ( .A1(dbg_uart_cmd[5]), .A2(dbg_uart_cmd[4]), .A3(
        dbg_uart_cmd[3]), .A4(n1518), .ZN(n2501) );
  inv0d0 U2254 ( .I(dbg_uart_cmd[2]), .ZN(n5960) );
  nd04d0 U2255 ( .A1(dbg_uart_cmd[0]), .A2(n1520), .A3(n2501), .A4(n5960), 
        .ZN(n1530) );
  oai21d1 U2256 ( .B1(dbg_uart_cmd[2]), .B2(dbg_uart_cmd[1]), .A(n2501), .ZN(
        n1519) );
  aoi211d1 U2257 ( .C1(dbg_uart_cmd[2]), .C2(dbg_uart_cmd[1]), .A(
        dbg_uart_cmd[0]), .B(n1519), .ZN(n2500) );
  nd02d0 U2258 ( .A1(n1520), .A2(n2500), .ZN(n1539) );
  oai211d1 U2259 ( .C1(n1521), .C2(n2504), .A(n1530), .B(n1539), .ZN(N6262) );
  nd02d0 U2260 ( .A1(n1524), .A2(n2482), .ZN(n1533) );
  inv0d0 U2261 ( .I(n1533), .ZN(n1528) );
  nr02d0 U2262 ( .A1(n1522), .A2(n5300), .ZN(n1523) );
  oan211d1 U2263 ( .C1(n1524), .C2(n5986), .B(n5489), .A(n1523), .ZN(n1534) );
  oai21d1 U2264 ( .B1(n1525), .B2(n5341), .A(n1534), .ZN(n1526) );
  oan211d1 U2265 ( .C1(n1528), .C2(n1527), .B(uartwishbonebridge_state[0]), 
        .A(n1526), .ZN(n1531) );
  nd02d0 U2266 ( .A1(uartwishbonebridge_state[0]), .A2(n1529), .ZN(n5968) );
  aon211d1 U2267 ( .C1(n1531), .C2(n5968), .B(n2504), .A(n1530), .ZN(N6263) );
  nr02d0 U2268 ( .A1(n1900), .A2(n1532), .ZN(n5297) );
  oai211d1 U2269 ( .C1(n5297), .C2(n1891), .A(n1534), .B(n1533), .ZN(n1537) );
  nr02d0 U2270 ( .A1(n5300), .A2(n1535), .ZN(n5320) );
  aoi22d1 U2271 ( .A1(uartwishbonebridge_state[2]), .A2(n1537), .B1(n5320), 
        .B2(n1536), .ZN(n1541) );
  inv0d0 U2272 ( .I(n1891), .ZN(n1898) );
  oai21d1 U2273 ( .B1(n1898), .B2(n1538), .A(uartwishbonebridge_state[0]), 
        .ZN(n1540) );
  aon211d1 U2274 ( .C1(n1541), .C2(n1540), .B(n2504), .A(n1539), .ZN(N6264) );
  nr02d0 U2275 ( .A1(litespi_state[0]), .A2(litespi_state[3]), .ZN(n1587) );
  oai21d1 U2276 ( .B1(litespi_state[2]), .B2(litespi_state[1]), .A(n1587), 
        .ZN(n1550) );
  nd12d0 U2277 ( .A1(n4684), .A2(n4685), .ZN(n1596) );
  nr04d0 U2278 ( .A1(mgmtsoc_litespisdrphycore_div[1]), .A2(
        mgmtsoc_litespisdrphycore_div[5]), .A3(
        mgmtsoc_litespisdrphycore_div[3]), .A4(
        mgmtsoc_litespisdrphycore_div[2]), .ZN(n1543) );
  nr04d0 U2279 ( .A1(mgmtsoc_litespisdrphycore_div[0]), .A2(
        mgmtsoc_litespisdrphycore_div[4]), .A3(
        mgmtsoc_litespisdrphycore_div[7]), .A4(
        mgmtsoc_litespisdrphycore_div[6]), .ZN(n1542) );
  nd02d0 U2280 ( .A1(n1543), .A2(n1542), .ZN(n5733) );
  nd02d0 U2281 ( .A1(n1544), .A2(litespiphy_state[1]), .ZN(n5734) );
  aoim21d1 U2282 ( .B1(mgmtsoc_litespisdrphycore_posedge_reg2), .B2(n5733), 
        .A(n5734), .ZN(n1599) );
  inv0d0 U2283 ( .I(n1599), .ZN(n1834) );
  nr02d0 U2284 ( .A1(litespi_tx_mux_sel), .A2(n1834), .ZN(n1552) );
  inv0d0 U2285 ( .I(n1552), .ZN(n1548) );
  nr03d0 U2286 ( .A1(mprj_we_o), .A2(n1545), .A3(n5050), .ZN(n1585) );
  inv0d0 U2287 ( .I(n1585), .ZN(n1930) );
  nd02d0 U2288 ( .A1(n1546), .A2(n1550), .ZN(n1606) );
  inv0d0 U2289 ( .I(n1551), .ZN(n4841) );
  nr02d0 U2290 ( .A1(n1606), .A2(n4841), .ZN(n4822) );
  inv0d0 U2291 ( .I(n4822), .ZN(n4843) );
  nr02d0 U2292 ( .A1(n1930), .A2(n4843), .ZN(n1547) );
  oan211d1 U2293 ( .C1(litespi_state[3]), .C2(n1548), .B(litespi_state[0]), 
        .A(n1547), .ZN(n1549) );
  oan211d1 U2294 ( .C1(n1550), .C2(n1596), .B(n1549), .A(n5492), .ZN(N6252) );
  nd02d0 U2295 ( .A1(n4822), .A2(n1930), .ZN(n1601) );
  aon211d1 U2296 ( .C1(litespi_state[0]), .C2(n1552), .B(litespi_state[3]), 
        .A(n1601), .ZN(n1591) );
  nr02d0 U2297 ( .A1(litespi_state[1]), .A2(n1551), .ZN(n1592) );
  aoi22d1 U2298 ( .A1(litespi_state[1]), .A2(n1591), .B1(n1592), .B2(n1552), 
        .ZN(n1589) );
  inv0d0 U2299 ( .I(mgmtsoc_litespimmap_spi_dummy_bits[4]), .ZN(n4816) );
  inv0d0 U2300 ( .I(mgmtsoc_litespimmap_spi_dummy_bits[5]), .ZN(n4817) );
  nd04d0 U2301 ( .A1(litespi_state[2]), .A2(n4816), .A3(n4817), .A4(n4815), 
        .ZN(n1554) );
  or04d0 U2302 ( .A1(mgmtsoc_litespimmap_spi_dummy_bits[0]), .A2(
        mgmtsoc_litespimmap_spi_dummy_bits[1]), .A3(
        mgmtsoc_litespimmap_spi_dummy_bits[2]), .A4(
        mgmtsoc_litespimmap_spi_dummy_bits[7]), .Z(n1553) );
  nr04d0 U2303 ( .A1(litespi_tx_mux_sel), .A2(n4684), .A3(n1554), .A4(n1553), 
        .ZN(n1586) );
  inv0d0 U2304 ( .I(mgmtsoc_litespimmap_spi_dummy_bits[6]), .ZN(n4818) );
  inv0d0 U2305 ( .I(mgmtsoc_litespimmap_burst_adr[0]), .ZN(n5609) );
  aoi22d1 U2306 ( .A1(n5611), .A2(n5609), .B1(mgmtsoc_litespimmap_burst_adr[0]), .B2(mprj_adr_o[2]), .ZN(n1584) );
  inv0d0 U2307 ( .I(mprj_adr_o[8]), .ZN(n5633) );
  oai22d1 U2308 ( .A1(n5625), .A2(mgmtsoc_litespimmap_burst_adr[4]), .B1(
        mgmtsoc_litespimmap_burst_adr[6]), .B2(n5633), .ZN(n1555) );
  aoi221d1 U2309 ( .B1(n5625), .B2(mgmtsoc_litespimmap_burst_adr[4]), .C1(
        n5633), .C2(mgmtsoc_litespimmap_burst_adr[6]), .A(n1555), .ZN(n1564)
         );
  oai22d1 U2310 ( .A1(n5629), .A2(mgmtsoc_litespimmap_burst_adr[5]), .B1(n5649), .B2(mgmtsoc_litespimmap_burst_adr[10]), .ZN(n1556) );
  aoi221d1 U2311 ( .B1(n5629), .B2(mgmtsoc_litespimmap_burst_adr[5]), .C1(
        mgmtsoc_litespimmap_burst_adr[10]), .C2(n5649), .A(n1556), .ZN(n1563)
         );
  inv0d0 U2312 ( .I(mgmtsoc_litespimmap_burst_adr[26]), .ZN(n1557) );
  nr04d0 U2313 ( .A1(mgmtsoc_litespimmap_burst_adr[27]), .A2(
        mgmtsoc_litespimmap_burst_adr[25]), .A3(
        mgmtsoc_litespimmap_burst_adr[24]), .A4(n1557), .ZN(n1562) );
  inv0d0 U2314 ( .I(mgmtsoc_litespimmap_burst_cs), .ZN(n1560) );
  aoi211d1 U2315 ( .C1(mgmtsoc_litespimmap_burst_adr[11]), .C2(n5653), .A(
        mgmtsoc_litespimmap_burst_adr[23]), .B(
        mgmtsoc_litespimmap_burst_adr[22]), .ZN(n1558) );
  oai21d1 U2316 ( .B1(mgmtsoc_litespimmap_burst_adr[11]), .B2(n5653), .A(n1558), .ZN(n1559) );
  oai22d1 U2317 ( .A1(n5670), .A2(mgmtsoc_litespimmap_burst_adr[15]), .B1(
        n5645), .B2(mgmtsoc_litespimmap_burst_adr[9]), .ZN(n1565) );
  aoi221d1 U2318 ( .B1(n5670), .B2(mgmtsoc_litespimmap_burst_adr[15]), .C1(
        mgmtsoc_litespimmap_burst_adr[9]), .C2(n5645), .A(n1565), .ZN(n1572)
         );
  oai22d1 U2319 ( .A1(n5674), .A2(mgmtsoc_litespimmap_burst_adr[16]), .B1(
        n5637), .B2(mgmtsoc_litespimmap_burst_adr[7]), .ZN(n1566) );
  aoi221d1 U2320 ( .B1(n5674), .B2(mgmtsoc_litespimmap_burst_adr[16]), .C1(
        mgmtsoc_litespimmap_burst_adr[7]), .C2(n5637), .A(n1566), .ZN(n1571)
         );
  inv0d0 U2321 ( .I(mprj_adr_o[20]), .ZN(n5682) );
  oai22d1 U2322 ( .A1(n5682), .A2(mgmtsoc_litespimmap_burst_adr[18]), .B1(
        n5614), .B2(mgmtsoc_litespimmap_burst_adr[1]), .ZN(n1567) );
  aoi221d1 U2323 ( .B1(n5682), .B2(mgmtsoc_litespimmap_burst_adr[18]), .C1(
        mgmtsoc_litespimmap_burst_adr[1]), .C2(n5614), .A(n1567), .ZN(n1570)
         );
  oai22d1 U2324 ( .A1(n5678), .A2(mgmtsoc_litespimmap_burst_adr[17]), .B1(
        mgmtsoc_litespimmap_burst_adr[2]), .B2(n5617), .ZN(n1568) );
  aoi221d1 U2325 ( .B1(n5678), .B2(mgmtsoc_litespimmap_burst_adr[17]), .C1(
        n5617), .C2(mgmtsoc_litespimmap_burst_adr[2]), .A(n1568), .ZN(n1569)
         );
  oai22d1 U2326 ( .A1(n5694), .A2(mgmtsoc_litespimmap_burst_adr[21]), .B1(
        n5657), .B2(mgmtsoc_litespimmap_burst_adr[12]), .ZN(n1573) );
  aoi221d1 U2327 ( .B1(n5694), .B2(mgmtsoc_litespimmap_burst_adr[21]), .C1(
        mgmtsoc_litespimmap_burst_adr[12]), .C2(n5657), .A(n1573), .ZN(n1580)
         );
  oai22d1 U2328 ( .A1(n5690), .A2(mgmtsoc_litespimmap_burst_adr[20]), .B1(
        n5661), .B2(mgmtsoc_litespimmap_burst_adr[13]), .ZN(n1574) );
  aoi221d1 U2329 ( .B1(n5690), .B2(mgmtsoc_litespimmap_burst_adr[20]), .C1(
        mgmtsoc_litespimmap_burst_adr[13]), .C2(n5661), .A(n1574), .ZN(n1579)
         );
  oai22d1 U2330 ( .A1(n5621), .A2(mgmtsoc_litespimmap_burst_adr[3]), .B1(n5641), .B2(mgmtsoc_litespimmap_burst_adr[8]), .ZN(n1575) );
  aoi221d1 U2331 ( .B1(n5621), .B2(mgmtsoc_litespimmap_burst_adr[3]), .C1(
        mgmtsoc_litespimmap_burst_adr[8]), .C2(n5641), .A(n1575), .ZN(n1578)
         );
  inv0d0 U2332 ( .I(mprj_adr_o[21]), .ZN(n5686) );
  oai22d1 U2333 ( .A1(n5666), .A2(mgmtsoc_litespimmap_burst_adr[14]), .B1(
        mgmtsoc_litespimmap_burst_adr[19]), .B2(n5686), .ZN(n1576) );
  aoi221d1 U2334 ( .B1(n5666), .B2(mgmtsoc_litespimmap_burst_adr[14]), .C1(
        n5686), .C2(mgmtsoc_litespimmap_burst_adr[19]), .A(n1576), .ZN(n1577)
         );
  nr04d0 U2335 ( .A1(n1584), .A2(n1583), .A3(n1582), .A4(n1581), .ZN(n1929) );
  an03d0 U2336 ( .A1(n1585), .A2(n1929), .A3(n4822), .Z(n1590) );
  aoi31d1 U2337 ( .B1(n1587), .B2(n1586), .B3(n4818), .A(n1590), .ZN(n1588) );
  aoi21d1 U2338 ( .B1(n1589), .B2(n1588), .A(n5100), .ZN(N6253) );
  oan211d1 U2339 ( .C1(n1592), .C2(n1591), .B(litespi_state[2]), .A(n1590), 
        .ZN(n1593) );
  oan211d1 U2340 ( .C1(n1834), .C2(n1594), .B(n1593), .A(sys_rst), .ZN(N6254)
         );
  nd02d0 U2341 ( .A1(litespi_state[2]), .A2(litespi_state[1]), .ZN(n4840) );
  aoi22d1 U2342 ( .A1(n1599), .A2(n1598), .B1(n1597), .B2(n1596), .ZN(n1600)
         );
  oan211d1 U2343 ( .C1(n1602), .C2(n1601), .B(n1600), .A(sys_rst), .ZN(N6255)
         );
  nr04d0 U2344 ( .A1(mgmtsoc_litespisdrphycore_sr_cnt[7]), .A2(
        mgmtsoc_litespisdrphycore_sr_cnt[6]), .A3(
        mgmtsoc_litespisdrphycore_sr_cnt[5]), .A4(
        mgmtsoc_litespisdrphycore_sr_cnt[4]), .ZN(n1604) );
  nr04d0 U2345 ( .A1(mgmtsoc_litespisdrphycore_sr_cnt[0]), .A2(
        mgmtsoc_litespisdrphycore_sr_cnt[1]), .A3(
        mgmtsoc_litespisdrphycore_sr_cnt[2]), .A4(
        mgmtsoc_litespisdrphycore_sr_cnt[3]), .ZN(n1603) );
  oan211d1 U2346 ( .C1(n4683), .C2(n4723), .B(
        \mgmtsoc_master_status_status[1] ), .A(n4685), .ZN(n4686) );
  aoi211d1 U2347 ( .C1(n4685), .C2(n1606), .A(n4686), .B(n4684), .ZN(n1608) );
  aoi211d1 U2348 ( .C1(n4857), .C2(n1609), .A(n5941), .B(n1608), .ZN(n1607) );
  aoi21d1 U2349 ( .B1(n1607), .B2(n1834), .A(n2516), .ZN(N6248) );
  inv0d0 U2350 ( .I(n1608), .ZN(n1610) );
  aoi31d1 U2351 ( .B1(n5734), .B2(n1610), .B3(n1609), .A(sys_rst), .ZN(N6249)
         );
  inv0d0 U2352 ( .I(n1611), .ZN(n1612) );
  oan211d1 U2353 ( .C1(csrbank9_cs0_w[16]), .C2(n1612), .B(csrbank9_cs0_w[0]), 
        .A(n5111), .ZN(N5589) );
  nr03d0 U2354 ( .A1(n5492), .A2(mgmtsoc_litespisdrphycore_clk), .A3(n1613), 
        .ZN(N5453) );
  inv0d0 U2355 ( .I(csrbank10_reload0_w[0]), .ZN(n4961) );
  nd02d0 U2356 ( .A1(csrbank10_en0_w), .A2(n5340), .ZN(n4954) );
  inv0d0 U2357 ( .I(n4954), .ZN(n1615) );
  nd02d1 U2358 ( .A1(n1614), .A2(n1615), .ZN(n1713) );
  buffd1 U2359 ( .I(n1713), .Z(n1702) );
  nd02d1 U2360 ( .A1(n4880), .A2(n1615), .ZN(n1712) );
  buffd1 U2361 ( .I(n1712), .Z(n1707) );
  inv0d0 U2362 ( .I(csrbank10_load0_w[0]), .ZN(n4999) );
  nd12d0 U2363 ( .A1(csrbank10_en0_w), .A2(n5301), .ZN(n1714) );
  buffd1 U2364 ( .I(n1714), .Z(n1703) );
  oai222d1 U2365 ( .A1(n4961), .A2(n1702), .B1(n1707), .B2(mgmtsoc_value[0]), 
        .C1(n4999), .C2(n1703), .ZN(N5400) );
  inv0d0 U2366 ( .I(csrbank10_load0_w[1]), .ZN(n5002) );
  inv0d0 U2367 ( .I(csrbank10_reload0_w[1]), .ZN(n4962) );
  inv0d0 U2368 ( .I(mgmtsoc_value[0]), .ZN(n4882) );
  aoim22d1 U2369 ( .A1(mgmtsoc_value[1]), .A2(n4882), .B1(n4882), .B2(
        mgmtsoc_value[1]), .Z(n1616) );
  inv0d0 U2370 ( .I(n1616), .ZN(n1617) );
  oai222d1 U2371 ( .A1(n1703), .A2(n5002), .B1(n1702), .B2(n4962), .C1(n1707), 
        .C2(n1617), .ZN(N5401) );
  inv0d0 U2372 ( .I(csrbank10_load0_w[2]), .ZN(n5003) );
  inv0d0 U2373 ( .I(csrbank10_reload0_w[2]), .ZN(n4963) );
  inv0d0 U2374 ( .I(mgmtsoc_value[2]), .ZN(n4887) );
  nr02d0 U2375 ( .A1(mgmtsoc_value[1]), .A2(mgmtsoc_value[0]), .ZN(n1618) );
  mi02d0 U2376 ( .I0(mgmtsoc_value[2]), .I1(n4887), .S(n1618), .ZN(n1619) );
  oai222d1 U2377 ( .A1(n1703), .A2(n5003), .B1(n1702), .B2(n4963), .C1(n1707), 
        .C2(n1619), .ZN(N5402) );
  inv0d0 U2378 ( .I(csrbank10_load0_w[3]), .ZN(n5005) );
  inv0d0 U2379 ( .I(csrbank10_reload0_w[3]), .ZN(n4964) );
  nr03d0 U2380 ( .A1(mgmtsoc_value[2]), .A2(mgmtsoc_value[1]), .A3(
        mgmtsoc_value[0]), .ZN(n1620) );
  aoim22d1 U2381 ( .A1(mgmtsoc_value[3]), .A2(n1620), .B1(n1620), .B2(
        mgmtsoc_value[3]), .Z(n1621) );
  inv0d0 U2382 ( .I(n1621), .ZN(n1622) );
  oai222d1 U2383 ( .A1(n1703), .A2(n5005), .B1(n1702), .B2(n4964), .C1(n1707), 
        .C2(n1622), .ZN(N5403) );
  inv0d0 U2384 ( .I(csrbank10_load0_w[4]), .ZN(n5007) );
  inv0d0 U2385 ( .I(csrbank10_reload0_w[4]), .ZN(n4965) );
  aoim22d1 U2386 ( .A1(mgmtsoc_value[4]), .A2(n1625), .B1(n1625), .B2(
        mgmtsoc_value[4]), .Z(n1623) );
  inv0d0 U2387 ( .I(n1623), .ZN(n1624) );
  oai222d1 U2388 ( .A1(n1703), .A2(n5007), .B1(n1702), .B2(n4965), .C1(n1707), 
        .C2(n1624), .ZN(N5404) );
  buffd1 U2389 ( .I(n1714), .Z(n1708) );
  inv0d0 U2390 ( .I(csrbank10_load0_w[5]), .ZN(n5009) );
  inv0d0 U2391 ( .I(csrbank10_reload0_w[5]), .ZN(n4966) );
  inv0d0 U2392 ( .I(mgmtsoc_value[5]), .ZN(n4893) );
  aoim22d1 U2393 ( .A1(n1628), .A2(n4893), .B1(n4893), .B2(n1628), .Z(n1626)
         );
  inv0d0 U2394 ( .I(n1626), .ZN(n1627) );
  oai222d1 U2395 ( .A1(n1708), .A2(n5009), .B1(n1713), .B2(n4966), .C1(n1712), 
        .C2(n1627), .ZN(N5405) );
  inv0d0 U2396 ( .I(csrbank10_load0_w[6]), .ZN(n5011) );
  inv0d0 U2397 ( .I(csrbank10_reload0_w[6]), .ZN(n4967) );
  nr02d0 U2398 ( .A1(n1628), .A2(mgmtsoc_value[5]), .ZN(n1631) );
  aoim22d1 U2399 ( .A1(mgmtsoc_value[6]), .A2(n1631), .B1(n1631), .B2(
        mgmtsoc_value[6]), .Z(n1629) );
  inv0d0 U2400 ( .I(n1629), .ZN(n1630) );
  oai222d1 U2401 ( .A1(n1708), .A2(n5011), .B1(n1713), .B2(n4967), .C1(n1712), 
        .C2(n1630), .ZN(N5406) );
  inv0d0 U2402 ( .I(csrbank10_load0_w[7]), .ZN(n5013) );
  inv0d0 U2403 ( .I(csrbank10_reload0_w[7]), .ZN(n4968) );
  nd12d0 U2404 ( .A1(mgmtsoc_value[6]), .A2(n1631), .ZN(n1634) );
  inv0d0 U2405 ( .I(mgmtsoc_value[7]), .ZN(n4897) );
  aoim22d1 U2406 ( .A1(n1634), .A2(n4897), .B1(n4897), .B2(n1634), .Z(n1632)
         );
  inv0d0 U2407 ( .I(n1632), .ZN(n1633) );
  oai222d1 U2408 ( .A1(n1708), .A2(n5013), .B1(n1702), .B2(n4968), .C1(n1712), 
        .C2(n1633), .ZN(N5407) );
  inv0d0 U2409 ( .I(csrbank10_load0_w[8]), .ZN(n5014) );
  inv0d0 U2410 ( .I(csrbank10_reload0_w[8]), .ZN(n4969) );
  nr02d0 U2411 ( .A1(n1634), .A2(mgmtsoc_value[7]), .ZN(n1637) );
  aoim22d1 U2412 ( .A1(mgmtsoc_value[8]), .A2(n1637), .B1(n1637), .B2(
        mgmtsoc_value[8]), .Z(n1635) );
  inv0d0 U2413 ( .I(n1635), .ZN(n1636) );
  oai222d1 U2414 ( .A1(n1708), .A2(n5014), .B1(n1713), .B2(n4969), .C1(n1712), 
        .C2(n1636), .ZN(N5408) );
  inv0d0 U2415 ( .I(csrbank10_load0_w[9]), .ZN(n5016) );
  inv0d0 U2416 ( .I(csrbank10_reload0_w[9]), .ZN(n4970) );
  nd12d0 U2417 ( .A1(mgmtsoc_value[8]), .A2(n1637), .ZN(n1641) );
  inv0d0 U2418 ( .I(n1641), .ZN(n1638) );
  aoim22d1 U2419 ( .A1(mgmtsoc_value[9]), .A2(n1638), .B1(n1638), .B2(
        mgmtsoc_value[9]), .Z(n1639) );
  inv0d0 U2420 ( .I(n1639), .ZN(n1640) );
  oai222d1 U2421 ( .A1(n1708), .A2(n5016), .B1(n1702), .B2(n4970), .C1(n1707), 
        .C2(n1640), .ZN(N5409) );
  inv0d0 U2422 ( .I(csrbank10_load0_w[10]), .ZN(n5018) );
  inv0d0 U2423 ( .I(csrbank10_reload0_w[10]), .ZN(n4971) );
  nr02d0 U2424 ( .A1(n1641), .A2(mgmtsoc_value[9]), .ZN(n1644) );
  aoim22d1 U2425 ( .A1(mgmtsoc_value[10]), .A2(n1644), .B1(n1644), .B2(
        mgmtsoc_value[10]), .Z(n1642) );
  inv0d0 U2426 ( .I(n1642), .ZN(n1643) );
  oai222d1 U2427 ( .A1(n1708), .A2(n5018), .B1(n1713), .B2(n4971), .C1(n1712), 
        .C2(n1643), .ZN(N5410) );
  inv0d0 U2428 ( .I(csrbank10_load0_w[11]), .ZN(n5020) );
  inv0d0 U2429 ( .I(csrbank10_reload0_w[11]), .ZN(n4972) );
  nd12d0 U2430 ( .A1(mgmtsoc_value[10]), .A2(n1644), .ZN(n1647) );
  inv0d0 U2431 ( .I(mgmtsoc_value[11]), .ZN(n4905) );
  aoim22d1 U2432 ( .A1(n1647), .A2(n4905), .B1(n4905), .B2(n1647), .Z(n1645)
         );
  inv0d0 U2433 ( .I(n1645), .ZN(n1646) );
  oai222d1 U2434 ( .A1(n1708), .A2(n5020), .B1(n1713), .B2(n4972), .C1(n1707), 
        .C2(n1646), .ZN(N5411) );
  inv0d0 U2435 ( .I(csrbank10_load0_w[12]), .ZN(n5021) );
  inv0d0 U2436 ( .I(csrbank10_reload0_w[12]), .ZN(n4973) );
  nr02d0 U2437 ( .A1(n1647), .A2(mgmtsoc_value[11]), .ZN(n1650) );
  aoim22d1 U2438 ( .A1(mgmtsoc_value[12]), .A2(n1650), .B1(n1650), .B2(
        mgmtsoc_value[12]), .Z(n1648) );
  inv0d0 U2439 ( .I(n1648), .ZN(n1649) );
  oai222d1 U2440 ( .A1(n1708), .A2(n5021), .B1(n1702), .B2(n4973), .C1(n1712), 
        .C2(n1649), .ZN(N5412) );
  inv0d0 U2441 ( .I(csrbank10_load0_w[13]), .ZN(n5023) );
  inv0d0 U2442 ( .I(csrbank10_reload0_w[13]), .ZN(n4974) );
  nd12d0 U2443 ( .A1(mgmtsoc_value[12]), .A2(n1650), .ZN(n1653) );
  inv0d0 U2444 ( .I(mgmtsoc_value[13]), .ZN(n4909) );
  aoim22d1 U2445 ( .A1(n1653), .A2(n4909), .B1(n4909), .B2(n1653), .Z(n1651)
         );
  inv0d0 U2446 ( .I(n1651), .ZN(n1652) );
  oai222d1 U2447 ( .A1(n1708), .A2(n5023), .B1(n1713), .B2(n4974), .C1(n1712), 
        .C2(n1652), .ZN(N5413) );
  inv0d0 U2448 ( .I(csrbank10_load0_w[14]), .ZN(n5025) );
  inv0d0 U2449 ( .I(csrbank10_reload0_w[14]), .ZN(n4975) );
  nr02d0 U2450 ( .A1(n1653), .A2(mgmtsoc_value[13]), .ZN(n1656) );
  aoim22d1 U2451 ( .A1(mgmtsoc_value[14]), .A2(n1656), .B1(n1656), .B2(
        mgmtsoc_value[14]), .Z(n1654) );
  inv0d0 U2452 ( .I(n1654), .ZN(n1655) );
  oai222d1 U2453 ( .A1(n1703), .A2(n5025), .B1(n1713), .B2(n4975), .C1(n1707), 
        .C2(n1655), .ZN(N5414) );
  inv0d0 U2454 ( .I(csrbank10_load0_w[15]), .ZN(n5027) );
  inv0d0 U2455 ( .I(csrbank10_reload0_w[15]), .ZN(n4976) );
  inv0d0 U2456 ( .I(mgmtsoc_value[15]), .ZN(n4913) );
  aoim22d1 U2457 ( .A1(n1657), .A2(n4913), .B1(n4913), .B2(n1657), .Z(n1658)
         );
  inv0d0 U2458 ( .I(n1658), .ZN(n1659) );
  oai222d1 U2459 ( .A1(n1703), .A2(n5027), .B1(n1702), .B2(n4976), .C1(n1707), 
        .C2(n1659), .ZN(N5415) );
  inv0d0 U2460 ( .I(csrbank10_load0_w[16]), .ZN(n5029) );
  inv0d0 U2461 ( .I(csrbank10_reload0_w[16]), .ZN(n4977) );
  inv0d0 U2462 ( .I(n1660), .ZN(n1663) );
  aoim22d1 U2463 ( .A1(mgmtsoc_value[16]), .A2(n1663), .B1(n1663), .B2(
        mgmtsoc_value[16]), .Z(n1661) );
  inv0d0 U2464 ( .I(n1661), .ZN(n1662) );
  oai222d1 U2465 ( .A1(n1708), .A2(n5029), .B1(n1713), .B2(n4977), .C1(n1712), 
        .C2(n1662), .ZN(N5416) );
  inv0d0 U2466 ( .I(csrbank10_load0_w[17]), .ZN(n5030) );
  inv0d0 U2467 ( .I(csrbank10_reload0_w[17]), .ZN(n4978) );
  nd12d0 U2468 ( .A1(mgmtsoc_value[16]), .A2(n1663), .ZN(n1666) );
  inv0d0 U2469 ( .I(mgmtsoc_value[17]), .ZN(n4917) );
  aoim22d1 U2470 ( .A1(n1666), .A2(n4917), .B1(n4917), .B2(n1666), .Z(n1664)
         );
  inv0d0 U2471 ( .I(n1664), .ZN(n1665) );
  oai222d1 U2472 ( .A1(n1708), .A2(n5030), .B1(n1702), .B2(n4978), .C1(n1712), 
        .C2(n1665), .ZN(N5417) );
  inv0d0 U2473 ( .I(csrbank10_load0_w[18]), .ZN(n5031) );
  inv0d0 U2474 ( .I(csrbank10_reload0_w[18]), .ZN(n4979) );
  nr02d0 U2475 ( .A1(n1666), .A2(mgmtsoc_value[17]), .ZN(n1669) );
  aoim22d1 U2476 ( .A1(mgmtsoc_value[18]), .A2(n1669), .B1(n1669), .B2(
        mgmtsoc_value[18]), .Z(n1667) );
  inv0d0 U2477 ( .I(n1667), .ZN(n1668) );
  oai222d1 U2478 ( .A1(n1703), .A2(n5031), .B1(n1702), .B2(n4979), .C1(n1712), 
        .C2(n1668), .ZN(N5418) );
  inv0d0 U2479 ( .I(csrbank10_load0_w[19]), .ZN(n5032) );
  inv0d0 U2480 ( .I(csrbank10_reload0_w[19]), .ZN(n4980) );
  nd12d0 U2481 ( .A1(mgmtsoc_value[18]), .A2(n1669), .ZN(n1672) );
  inv0d0 U2482 ( .I(mgmtsoc_value[19]), .ZN(n4921) );
  aoim22d1 U2483 ( .A1(n1672), .A2(n4921), .B1(n4921), .B2(n1672), .Z(n1670)
         );
  inv0d0 U2484 ( .I(n1670), .ZN(n1671) );
  oai222d1 U2485 ( .A1(n1703), .A2(n5032), .B1(n1702), .B2(n4980), .C1(n1712), 
        .C2(n1671), .ZN(N5419) );
  inv0d0 U2486 ( .I(csrbank10_load0_w[20]), .ZN(n5033) );
  inv0d0 U2487 ( .I(csrbank10_reload0_w[20]), .ZN(n4981) );
  nr02d0 U2488 ( .A1(n1672), .A2(mgmtsoc_value[19]), .ZN(n1675) );
  aoim22d1 U2489 ( .A1(mgmtsoc_value[20]), .A2(n1675), .B1(n1675), .B2(
        mgmtsoc_value[20]), .Z(n1673) );
  inv0d0 U2490 ( .I(n1673), .ZN(n1674) );
  oai222d1 U2491 ( .A1(n1703), .A2(n5033), .B1(n1713), .B2(n4981), .C1(n1707), 
        .C2(n1674), .ZN(N5420) );
  inv0d0 U2492 ( .I(csrbank10_load0_w[21]), .ZN(n5034) );
  inv0d0 U2493 ( .I(csrbank10_reload0_w[21]), .ZN(n4982) );
  nd12d0 U2494 ( .A1(mgmtsoc_value[20]), .A2(n1675), .ZN(n1678) );
  inv0d0 U2495 ( .I(mgmtsoc_value[21]), .ZN(n4925) );
  aoim22d1 U2496 ( .A1(n1678), .A2(n4925), .B1(n4925), .B2(n1678), .Z(n1676)
         );
  inv0d0 U2497 ( .I(n1676), .ZN(n1677) );
  oai222d1 U2498 ( .A1(n1708), .A2(n5034), .B1(n1702), .B2(n4982), .C1(n1712), 
        .C2(n1677), .ZN(N5421) );
  inv0d0 U2499 ( .I(csrbank10_load0_w[22]), .ZN(n5035) );
  inv0d0 U2500 ( .I(csrbank10_reload0_w[22]), .ZN(n4983) );
  nr02d0 U2501 ( .A1(n1678), .A2(mgmtsoc_value[21]), .ZN(n1681) );
  aoim22d1 U2502 ( .A1(mgmtsoc_value[22]), .A2(n1681), .B1(n1681), .B2(
        mgmtsoc_value[22]), .Z(n1679) );
  inv0d0 U2503 ( .I(n1679), .ZN(n1680) );
  oai222d1 U2504 ( .A1(n1703), .A2(n5035), .B1(n1713), .B2(n4983), .C1(n1707), 
        .C2(n1680), .ZN(N5422) );
  inv0d0 U2505 ( .I(csrbank10_load0_w[23]), .ZN(n5036) );
  inv0d0 U2506 ( .I(csrbank10_reload0_w[23]), .ZN(n4984) );
  inv0d0 U2507 ( .I(mgmtsoc_value[23]), .ZN(n4929) );
  aoim22d1 U2508 ( .A1(n1684), .A2(n4929), .B1(n4929), .B2(n1684), .Z(n1682)
         );
  inv0d0 U2509 ( .I(n1682), .ZN(n1683) );
  oai222d1 U2510 ( .A1(n1703), .A2(n5036), .B1(n1702), .B2(n4984), .C1(n1707), 
        .C2(n1683), .ZN(N5423) );
  inv0d0 U2511 ( .I(csrbank10_load0_w[24]), .ZN(n5037) );
  inv0d0 U2512 ( .I(csrbank10_reload0_w[24]), .ZN(n4985) );
  nr02d0 U2513 ( .A1(n1684), .A2(mgmtsoc_value[23]), .ZN(n1687) );
  aoim22d1 U2514 ( .A1(mgmtsoc_value[24]), .A2(n1687), .B1(n1687), .B2(
        mgmtsoc_value[24]), .Z(n1685) );
  inv0d0 U2515 ( .I(n1685), .ZN(n1686) );
  oai222d1 U2516 ( .A1(n1703), .A2(n5037), .B1(n1713), .B2(n4985), .C1(n1707), 
        .C2(n1686), .ZN(N5424) );
  inv0d0 U2517 ( .I(csrbank10_load0_w[25]), .ZN(n5039) );
  inv0d0 U2518 ( .I(csrbank10_reload0_w[25]), .ZN(n4986) );
  nd12d0 U2519 ( .A1(mgmtsoc_value[24]), .A2(n1687), .ZN(n1690) );
  inv0d0 U2520 ( .I(mgmtsoc_value[25]), .ZN(n4933) );
  aoim22d1 U2521 ( .A1(n1690), .A2(n4933), .B1(n4933), .B2(n1690), .Z(n1688)
         );
  inv0d0 U2522 ( .I(n1688), .ZN(n1689) );
  oai222d1 U2523 ( .A1(n1708), .A2(n5039), .B1(n1713), .B2(n4986), .C1(n1707), 
        .C2(n1689), .ZN(N5425) );
  inv0d0 U2524 ( .I(csrbank10_load0_w[26]), .ZN(n5040) );
  inv0d0 U2525 ( .I(csrbank10_reload0_w[26]), .ZN(n4988) );
  nr02d0 U2526 ( .A1(n1690), .A2(mgmtsoc_value[25]), .ZN(n1693) );
  aoim22d1 U2527 ( .A1(mgmtsoc_value[26]), .A2(n1693), .B1(n1693), .B2(
        mgmtsoc_value[26]), .Z(n1691) );
  inv0d0 U2528 ( .I(n1691), .ZN(n1692) );
  oai222d1 U2529 ( .A1(n1703), .A2(n5040), .B1(n1713), .B2(n4988), .C1(n1707), 
        .C2(n1692), .ZN(N5426) );
  inv0d0 U2530 ( .I(csrbank10_load0_w[27]), .ZN(n5041) );
  inv0d0 U2531 ( .I(csrbank10_reload0_w[27]), .ZN(n4989) );
  inv0d0 U2532 ( .I(mgmtsoc_value[27]), .ZN(n4938) );
  aoim22d1 U2533 ( .A1(n1696), .A2(n4938), .B1(n4938), .B2(n1696), .Z(n1694)
         );
  inv0d0 U2534 ( .I(n1694), .ZN(n1695) );
  oai222d1 U2535 ( .A1(n1708), .A2(n5041), .B1(n1702), .B2(n4989), .C1(n1707), 
        .C2(n1695), .ZN(N5427) );
  inv0d0 U2536 ( .I(csrbank10_load0_w[28]), .ZN(n5042) );
  inv0d0 U2537 ( .I(csrbank10_reload0_w[28]), .ZN(n4990) );
  nr02d0 U2538 ( .A1(n1696), .A2(mgmtsoc_value[27]), .ZN(n1699) );
  aoim22d1 U2539 ( .A1(mgmtsoc_value[28]), .A2(n1699), .B1(n1699), .B2(
        mgmtsoc_value[28]), .Z(n1697) );
  inv0d0 U2540 ( .I(n1697), .ZN(n1698) );
  oai222d1 U2541 ( .A1(n1714), .A2(n5042), .B1(n1702), .B2(n4990), .C1(n1712), 
        .C2(n1698), .ZN(N5428) );
  inv0d0 U2542 ( .I(csrbank10_load0_w[29]), .ZN(n5043) );
  inv0d0 U2543 ( .I(csrbank10_reload0_w[29]), .ZN(n4992) );
  inv0d0 U2544 ( .I(mgmtsoc_value[29]), .ZN(n4942) );
  aoim22d1 U2545 ( .A1(n1704), .A2(n4942), .B1(n4942), .B2(n1704), .Z(n1700)
         );
  inv0d0 U2546 ( .I(n1700), .ZN(n1701) );
  oai222d1 U2547 ( .A1(n1703), .A2(n5043), .B1(n1702), .B2(n4992), .C1(n1712), 
        .C2(n1701), .ZN(N5429) );
  inv0d0 U2548 ( .I(csrbank10_load0_w[30]), .ZN(n5044) );
  inv0d0 U2549 ( .I(csrbank10_reload0_w[30]), .ZN(n4993) );
  nr02d0 U2550 ( .A1(n1704), .A2(mgmtsoc_value[29]), .ZN(n1709) );
  aoim22d1 U2551 ( .A1(mgmtsoc_value[30]), .A2(n1709), .B1(n1709), .B2(
        mgmtsoc_value[30]), .Z(n1705) );
  inv0d0 U2552 ( .I(n1705), .ZN(n1706) );
  oai222d1 U2553 ( .A1(n1708), .A2(n5044), .B1(n1713), .B2(n4993), .C1(n1707), 
        .C2(n1706), .ZN(N5430) );
  inv0d0 U2554 ( .I(csrbank10_load0_w[31]), .ZN(n5047) );
  inv0d0 U2555 ( .I(csrbank10_reload0_w[31]), .ZN(n4995) );
  inv0d0 U2556 ( .I(n1709), .ZN(n1710) );
  oai21d1 U2557 ( .B1(mgmtsoc_value[30]), .B2(n1710), .A(mgmtsoc_value[31]), 
        .ZN(n1711) );
  oai222d1 U2558 ( .A1(n1714), .A2(n5047), .B1(n1713), .B2(n4995), .C1(n1712), 
        .C2(n1711), .ZN(N5431) );
  ah01d1 U2559 ( .A(n1715), .B(dbg_uart_rx_phase[31]), .CO(n1277), .S(n1716)
         );
  aoim21d1 U2560 ( .B1(n1716), .B2(n2874), .A(n5492), .ZN(N5077) );
  inv0d0 U2561 ( .I(dbg_uart_tx_phase[0]), .ZN(n1717) );
  nr02d0 U2562 ( .A1(n5492), .A2(uartwishbonebridge_rs232phytx_state), .ZN(
        n2508) );
  inv0d1 U2563 ( .I(n2508), .ZN(n5988) );
  oaim21d1 U2564 ( .B1(n1717), .B2(n5956), .A(n5988), .ZN(N5014) );
  aoim22d1 U2565 ( .A1(dbg_uart_tx_phase[1]), .A2(n1717), .B1(n1717), .B2(
        dbg_uart_tx_phase[1]), .Z(n1718) );
  oaim21d1 U2566 ( .B1(n1718), .B2(n5301), .A(n5988), .ZN(N5015) );
  mx02d1 U2567 ( .I0(dbg_uart_tx_phase[2]), .I1(n1720), .S(n1719), .Z(n1721)
         );
  oaim21d1 U2568 ( .B1(n1721), .B2(n5956), .A(n5988), .ZN(N5016) );
  inv0d0 U2569 ( .I(n1722), .ZN(n1723) );
  aoim22d1 U2570 ( .A1(dbg_uart_tx_phase[7]), .A2(n1723), .B1(n1723), .B2(
        dbg_uart_tx_phase[7]), .Z(n1724) );
  oaim21d1 U2571 ( .B1(n1724), .B2(n5956), .A(n5988), .ZN(N5021) );
  mx02d1 U2572 ( .I0(dbg_uart_tx_phase[8]), .I1(n1726), .S(n1725), .Z(n1727)
         );
  oaim21d1 U2573 ( .B1(n1727), .B2(n5956), .A(n5988), .ZN(N5022) );
  inv0d0 U2574 ( .I(n1730), .ZN(n1728) );
  aoim22d1 U2575 ( .A1(dbg_uart_tx_phase[11]), .A2(n1728), .B1(n1728), .B2(
        dbg_uart_tx_phase[11]), .Z(n1729) );
  oaim21d1 U2576 ( .B1(n1729), .B2(n5340), .A(n5988), .ZN(N5025) );
  inv0d0 U2577 ( .I(dbg_uart_tx_phase[12]), .ZN(n1732) );
  nr02d0 U2578 ( .A1(dbg_uart_tx_phase[11]), .A2(n1730), .ZN(n1731) );
  mx02d1 U2579 ( .I0(dbg_uart_tx_phase[12]), .I1(n1732), .S(n1731), .Z(n1733)
         );
  oaim21d1 U2580 ( .B1(n1733), .B2(n5956), .A(n5988), .ZN(N5026) );
  aoim22d1 U2581 ( .A1(dbg_uart_tx_phase[13]), .A2(n1734), .B1(n1734), .B2(
        dbg_uart_tx_phase[13]), .Z(n1735) );
  oaim21d1 U2582 ( .B1(n1735), .B2(n5301), .A(n5988), .ZN(N5027) );
  inv0d0 U2583 ( .I(n1736), .ZN(n1737) );
  aoim22d1 U2584 ( .A1(dbg_uart_tx_phase[14]), .A2(n1737), .B1(n1737), .B2(
        dbg_uart_tx_phase[14]), .Z(n1738) );
  oaim21d1 U2585 ( .B1(n1738), .B2(n5956), .A(n5988), .ZN(N5028) );
  mx02d1 U2586 ( .I0(dbg_uart_tx_phase[15]), .I1(n1740), .S(n1739), .Z(n1741)
         );
  oaim21d1 U2587 ( .B1(n1741), .B2(n4881), .A(n5988), .ZN(N5029) );
  aoi22d1 U2588 ( .A1(dbg_uart_tx_phase[17]), .A2(n1744), .B1(n1743), .B2(
        n1742), .ZN(n1745) );
  oaim21d1 U2589 ( .B1(n1745), .B2(n5340), .A(n5988), .ZN(N5031) );
  inv0d0 U2590 ( .I(n1751), .ZN(n1746) );
  aoim22d1 U2591 ( .A1(dbg_uart_tx_phase[20]), .A2(n1746), .B1(n1746), .B2(
        dbg_uart_tx_phase[20]), .Z(n1747) );
  oaim21d1 U2592 ( .B1(n1747), .B2(n5340), .A(n5988), .ZN(N5034) );
  inv0d0 U2593 ( .I(dbg_uart_tx_phase[21]), .ZN(n1749) );
  mx02d1 U2594 ( .I0(dbg_uart_tx_phase[21]), .I1(n1749), .S(n1748), .Z(n1750)
         );
  oaim21d1 U2595 ( .B1(n1750), .B2(n5340), .A(n5988), .ZN(N5035) );
  inv0d0 U2596 ( .I(dbg_uart_tx_phase[22]), .ZN(n1753) );
  nr03d0 U2597 ( .A1(dbg_uart_tx_phase[21]), .A2(dbg_uart_tx_phase[20]), .A3(
        n1751), .ZN(n1752) );
  mx02d1 U2598 ( .I0(dbg_uart_tx_phase[22]), .I1(n1753), .S(n1752), .Z(n1754)
         );
  oaim21d1 U2599 ( .B1(n1754), .B2(n5956), .A(n5988), .ZN(N5036) );
  mx02d1 U2600 ( .I0(dbg_uart_tx_phase[23]), .I1(n1756), .S(n1755), .Z(n1757)
         );
  oaim21d1 U2601 ( .B1(n1757), .B2(n4881), .A(n5988), .ZN(N5037) );
  aoi22d1 U2602 ( .A1(dbg_uart_tx_phase[25]), .A2(n1760), .B1(n1759), .B2(
        n1758), .ZN(n1761) );
  oaim21d1 U2603 ( .B1(n1761), .B2(n4881), .A(n5988), .ZN(N5039) );
  inv0d0 U2604 ( .I(csrbank18_edge0_w), .ZN(n1771) );
  nr02d0 U2605 ( .A1(n1783), .A2(n1762), .ZN(n1763) );
  aoi22d1 U2606 ( .A1(n2476), .A2(csrbank18_in_w), .B1(gpioin5_i01), .B2(n1763), .ZN(n1767) );
  nd13d1 U2607 ( .A1(n1934), .A2(n1765), .A3(n1764), .ZN(n1766) );
  oai211d1 U2608 ( .C1(n1847), .C2(n1768), .A(n1767), .B(n1766), .ZN(n1769) );
  aoi31d1 U2609 ( .B1(n1903), .B2(n1902), .B3(gpioin5_i02), .A(n1769), .ZN(
        n1770) );
  oan211d1 U2610 ( .C1(n1846), .C2(n1771), .B(n1770), .A(n1937), .ZN(N4982) );
  aoi22d1 U2611 ( .A1(n4998), .A2(csrbank16_in_w), .B1(n1839), .B2(gpioin3_i01), .ZN(n1775) );
  aoim22d1 U2612 ( .A1(n4952), .A2(csrbank16_edge0_w), .B1(n2451), .B2(n1949), 
        .Z(n1774) );
  aoi22d1 U2613 ( .A1(n1902), .A2(gpioin3_i02), .B1(n2457), .B2(
        csrbank16_mode0_w), .ZN(n1773) );
  nd02d0 U2614 ( .A1(n1903), .A2(n1912), .ZN(n1772) );
  aoi31d1 U2615 ( .B1(n1775), .B2(n1774), .B3(n1773), .A(n1772), .ZN(N4918) );
  oai21d1 U2616 ( .B1(csrbank15_mode0_w), .B2(n2451), .A(n2454), .ZN(n1776) );
  aoi22d1 U2617 ( .A1(n2457), .A2(csrbank15_mode0_w), .B1(csrbank15_edge0_w), 
        .B2(n1776), .ZN(n1778) );
  aoi22d1 U2618 ( .A1(n1902), .A2(gpioin2_i02), .B1(n1839), .B2(gpioin2_i01), 
        .ZN(n1777) );
  aoi211d1 U2619 ( .C1(n1778), .C2(n1777), .A(n1959), .B(n1783), .ZN(N4886) );
  oai21d1 U2620 ( .B1(csrbank14_mode0_w), .B2(n2451), .A(n2454), .ZN(n1779) );
  aoi22d1 U2621 ( .A1(n2457), .A2(csrbank14_mode0_w), .B1(csrbank14_edge0_w), 
        .B2(n1779), .ZN(n1781) );
  aoi22d1 U2622 ( .A1(n1902), .A2(gpioin1_i02), .B1(n1839), .B2(gpioin1_i01), 
        .ZN(n1780) );
  aoi211d1 U2623 ( .C1(n1781), .C2(n1780), .A(n1966), .B(n1783), .ZN(N4854) );
  oai21d1 U2624 ( .B1(csrbank13_mode0_w), .B2(n2451), .A(n2454), .ZN(n1782) );
  aoi22d1 U2625 ( .A1(n2457), .A2(csrbank13_mode0_w), .B1(csrbank13_edge0_w), 
        .B2(n1782), .ZN(n1785) );
  aoi22d1 U2626 ( .A1(n1902), .A2(gpioin0_i02), .B1(n1839), .B2(gpioin0_i01), 
        .ZN(n1784) );
  aoi211d1 U2627 ( .C1(n1785), .C2(n1784), .A(n1973), .B(n1783), .ZN(N4822) );
  inv0d0 U2628 ( .I(uart_phy_tx_sink_valid), .ZN(n2666) );
  aoi22d1 U2629 ( .A1(csrbank11_ev_enable0_w[0]), .A2(n1902), .B1(n1806), .B2(
        n2666), .ZN(n1790) );
  aoi22d1 U2630 ( .A1(n4998), .A2(uart_rx_fifo_fifo_out_payload_data[0]), .B1(
        n1839), .B2(uart_pending_status[0]), .ZN(n1789) );
  nr04d0 U2631 ( .A1(uart_rx_fifo_level0[3]), .A2(uart_rx_fifo_level0[2]), 
        .A3(uart_rx_fifo_level0[1]), .A4(uart_rx_fifo_level0[0]), .ZN(n2550)
         );
  nd02d0 U2632 ( .A1(uart_rx_fifo_level0[4]), .A2(n2550), .ZN(n2518) );
  oai22d1 U2633 ( .A1(\uart_status_status[1] ), .A2(n2454), .B1(n1786), .B2(
        n2518), .ZN(n1787) );
  aoi221d1 U2634 ( .B1(n2457), .B2(n2664), .C1(n1838), .C2(n2556), .A(n1787), 
        .ZN(n1788) );
  inv0d0 U2635 ( .I(n2655), .ZN(n2648) );
  nd02d0 U2636 ( .A1(n1903), .A2(n2648), .ZN(n1791) );
  aoi31d1 U2637 ( .B1(n1790), .B2(n1789), .B3(n1788), .A(n1791), .ZN(N4772) );
  aoi22d1 U2638 ( .A1(n1838), .A2(\uart_status_status[1] ), .B1(n1902), .B2(
        csrbank11_ev_enable0_w[1]), .ZN(n1793) );
  aoi22d1 U2639 ( .A1(n4998), .A2(uart_rx_fifo_fifo_out_payload_data[1]), .B1(
        n1839), .B2(uart_pending_status[1]), .ZN(n1792) );
  aoi21d1 U2640 ( .B1(n1793), .B2(n1792), .A(n1791), .ZN(N4773) );
  nd02d1 U2641 ( .A1(n1839), .A2(n1794), .ZN(n1797) );
  buffd1 U2642 ( .I(n1797), .Z(n1798) );
  inv0d0 U2643 ( .I(csrbank10_value_w[1]), .ZN(n4884) );
  nd02d1 U2644 ( .A1(n2457), .A2(n1794), .ZN(n1795) );
  buffd1 U2645 ( .I(n1795), .Z(n4958) );
  nd12d1 U2646 ( .A1(n4960), .A2(n2476), .ZN(n1796) );
  buffd1 U2647 ( .I(n1796), .Z(n1799) );
  oai222d1 U2648 ( .A1(n1798), .A2(n4884), .B1(n4962), .B2(n4958), .C1(n5002), 
        .C2(n1799), .ZN(N4695) );
  inv0d0 U2649 ( .I(csrbank10_value_w[2]), .ZN(n4886) );
  oai222d1 U2650 ( .A1(n5003), .A2(n1799), .B1(n4963), .B2(n1795), .C1(n4886), 
        .C2(n1797), .ZN(N4696) );
  inv0d0 U2651 ( .I(csrbank10_value_w[3]), .ZN(n4888) );
  oai222d1 U2652 ( .A1(n5005), .A2(n1799), .B1(n4964), .B2(n4958), .C1(n1798), 
        .C2(n4888), .ZN(N4697) );
  inv0d0 U2653 ( .I(csrbank10_value_w[4]), .ZN(n4890) );
  oai222d1 U2654 ( .A1(n5007), .A2(n1799), .B1(n4965), .B2(n4958), .C1(n1798), 
        .C2(n4890), .ZN(N4698) );
  inv0d0 U2655 ( .I(csrbank10_value_w[5]), .ZN(n4892) );
  oai222d1 U2656 ( .A1(n5009), .A2(n1799), .B1(n4966), .B2(n4958), .C1(n1798), 
        .C2(n4892), .ZN(N4699) );
  inv0d0 U2657 ( .I(csrbank10_value_w[6]), .ZN(n4894) );
  oai222d1 U2658 ( .A1(n5011), .A2(n1799), .B1(n4967), .B2(n1795), .C1(n4894), 
        .C2(n1797), .ZN(N4700) );
  inv0d0 U2659 ( .I(csrbank10_value_w[7]), .ZN(n4896) );
  oai222d1 U2660 ( .A1(n5013), .A2(n1799), .B1(n4968), .B2(n1795), .C1(n1798), 
        .C2(n4896), .ZN(N4701) );
  inv0d0 U2661 ( .I(csrbank10_value_w[8]), .ZN(n4898) );
  oai222d1 U2662 ( .A1(n5014), .A2(n1799), .B1(n4969), .B2(n1795), .C1(n4898), 
        .C2(n1797), .ZN(N4702) );
  inv0d0 U2663 ( .I(csrbank10_value_w[9]), .ZN(n4900) );
  oai222d1 U2664 ( .A1(n5016), .A2(n1799), .B1(n4970), .B2(n4958), .C1(n4900), 
        .C2(n1797), .ZN(N4703) );
  inv0d0 U2665 ( .I(csrbank10_value_w[10]), .ZN(n4902) );
  oai222d1 U2666 ( .A1(n5018), .A2(n1796), .B1(n4971), .B2(n4958), .C1(n1798), 
        .C2(n4902), .ZN(N4704) );
  inv0d0 U2667 ( .I(csrbank10_value_w[11]), .ZN(n4904) );
  oai222d1 U2668 ( .A1(n5020), .A2(n1799), .B1(n4972), .B2(n4958), .C1(n4904), 
        .C2(n1797), .ZN(N4705) );
  inv0d0 U2669 ( .I(csrbank10_value_w[12]), .ZN(n4906) );
  oai222d1 U2670 ( .A1(n5021), .A2(n1799), .B1(n4973), .B2(n4958), .C1(n4906), 
        .C2(n1797), .ZN(N4706) );
  inv0d0 U2671 ( .I(csrbank10_value_w[13]), .ZN(n4908) );
  oai222d1 U2672 ( .A1(n5023), .A2(n1796), .B1(n4974), .B2(n1795), .C1(n4908), 
        .C2(n1798), .ZN(N4707) );
  inv0d0 U2673 ( .I(csrbank10_value_w[14]), .ZN(n4910) );
  oai222d1 U2674 ( .A1(n5025), .A2(n1796), .B1(n4975), .B2(n4958), .C1(n1798), 
        .C2(n4910), .ZN(N4708) );
  inv0d0 U2675 ( .I(csrbank10_value_w[15]), .ZN(n4912) );
  oai222d1 U2676 ( .A1(n5027), .A2(n1796), .B1(n4976), .B2(n1795), .C1(n4912), 
        .C2(n1797), .ZN(N4709) );
  inv0d0 U2677 ( .I(csrbank10_value_w[16]), .ZN(n4914) );
  oai222d1 U2678 ( .A1(n5029), .A2(n1796), .B1(n4977), .B2(n1795), .C1(n4914), 
        .C2(n1798), .ZN(N4710) );
  inv0d0 U2679 ( .I(csrbank10_value_w[17]), .ZN(n4916) );
  oai222d1 U2680 ( .A1(n5030), .A2(n1799), .B1(n4978), .B2(n1795), .C1(n4916), 
        .C2(n1797), .ZN(N4711) );
  inv0d0 U2681 ( .I(csrbank10_value_w[18]), .ZN(n4918) );
  oai222d1 U2682 ( .A1(n5031), .A2(n1796), .B1(n4979), .B2(n4958), .C1(n4918), 
        .C2(n1797), .ZN(N4712) );
  inv0d0 U2683 ( .I(csrbank10_value_w[19]), .ZN(n4920) );
  oai222d1 U2684 ( .A1(n5032), .A2(n1799), .B1(n4980), .B2(n1795), .C1(n4920), 
        .C2(n1798), .ZN(N4713) );
  inv0d0 U2685 ( .I(csrbank10_value_w[20]), .ZN(n4922) );
  oai222d1 U2686 ( .A1(n5033), .A2(n1796), .B1(n4981), .B2(n1795), .C1(n1798), 
        .C2(n4922), .ZN(N4714) );
  inv0d0 U2687 ( .I(csrbank10_value_w[21]), .ZN(n4924) );
  oai222d1 U2688 ( .A1(n5034), .A2(n1796), .B1(n4982), .B2(n4958), .C1(n1797), 
        .C2(n4924), .ZN(N4715) );
  inv0d0 U2689 ( .I(csrbank10_value_w[22]), .ZN(n4926) );
  oai222d1 U2690 ( .A1(n5035), .A2(n1799), .B1(n4983), .B2(n4958), .C1(n4926), 
        .C2(n1798), .ZN(N4716) );
  inv0d0 U2691 ( .I(csrbank10_value_w[23]), .ZN(n4928) );
  oai222d1 U2692 ( .A1(n5036), .A2(n1796), .B1(n4984), .B2(n1795), .C1(n4928), 
        .C2(n1797), .ZN(N4717) );
  inv0d0 U2693 ( .I(csrbank10_value_w[24]), .ZN(n4930) );
  oai222d1 U2694 ( .A1(n5037), .A2(n1796), .B1(n4985), .B2(n1795), .C1(n1798), 
        .C2(n4930), .ZN(N4718) );
  inv0d0 U2695 ( .I(csrbank10_value_w[25]), .ZN(n4932) );
  oai222d1 U2696 ( .A1(n5039), .A2(n1796), .B1(n4986), .B2(n1795), .C1(n4932), 
        .C2(n1797), .ZN(N4719) );
  inv0d0 U2697 ( .I(csrbank10_value_w[26]), .ZN(n4935) );
  oai222d1 U2698 ( .A1(n5040), .A2(n1796), .B1(n4988), .B2(n1795), .C1(n4935), 
        .C2(n1798), .ZN(N4720) );
  inv0d0 U2699 ( .I(csrbank10_value_w[27]), .ZN(n4937) );
  oai222d1 U2700 ( .A1(n5041), .A2(n1796), .B1(n4989), .B2(n1795), .C1(n4937), 
        .C2(n1797), .ZN(N4721) );
  inv0d0 U2701 ( .I(csrbank10_value_w[28]), .ZN(n4939) );
  oai222d1 U2702 ( .A1(n5042), .A2(n1799), .B1(n4990), .B2(n4958), .C1(n1798), 
        .C2(n4939), .ZN(N4722) );
  inv0d0 U2703 ( .I(csrbank10_value_w[29]), .ZN(n4941) );
  oai222d1 U2704 ( .A1(n5043), .A2(n1796), .B1(n4992), .B2(n4958), .C1(n1798), 
        .C2(n4941), .ZN(N4723) );
  inv0d0 U2705 ( .I(csrbank10_value_w[30]), .ZN(n4943) );
  oai222d1 U2706 ( .A1(n5044), .A2(n1799), .B1(n4993), .B2(n4958), .C1(n4943), 
        .C2(n1797), .ZN(N4724) );
  inv0d0 U2707 ( .I(csrbank10_value_w[31]), .ZN(n4947) );
  oai222d1 U2708 ( .A1(n5047), .A2(n1799), .B1(n4995), .B2(n4958), .C1(n4947), 
        .C2(n1798), .ZN(N4725) );
  aoi211d1 U2709 ( .C1(csrbank9_control0_w[0]), .C2(spi_master_control_re), 
        .A(spimaster_state[1]), .B(spimaster_state[0]), .ZN(n1800) );
  aoi22d1 U2710 ( .A1(n1838), .A2(spi_master_miso_status[0]), .B1(n2457), .B2(
        n1800), .ZN(n1804) );
  aoi22d1 U2711 ( .A1(n1806), .A2(spi_master_clk_divider0[0]), .B1(n4952), 
        .B2(spi_master_mosi[0]), .ZN(n1803) );
  aor22d1 U2712 ( .A1(n4998), .A2(csrbank9_control0_w[0]), .B1(n1839), .B2(
        csrbank9_cs0_w[0]), .Z(n1801) );
  aoi21d1 U2713 ( .B1(n1902), .B2(spi_master_loopback), .A(n1801), .ZN(n1802)
         );
  aoi31d1 U2714 ( .B1(n1804), .B2(n1803), .B3(n1802), .A(n1807), .ZN(N4585) );
  nd02d1 U2715 ( .A1(n1806), .A2(n1805), .ZN(n1827) );
  inv0d0 U2716 ( .I(spi_master_clk_divider0[1]), .ZN(n3064) );
  aoi22d1 U2717 ( .A1(n4579), .A2(csrbank9_cs0_w[1]), .B1(
        spi_master_miso_status[1]), .B2(n1822), .ZN(n1809) );
  nr02d0 U2718 ( .A1(n1807), .A2(n2454), .ZN(n1818) );
  aoi22d1 U2719 ( .A1(spi_master_mosi[1]), .A2(n1818), .B1(n1821), .B2(
        csrbank9_control0_w[1]), .ZN(n1808) );
  oai211d1 U2720 ( .C1(n1827), .C2(n3064), .A(n1809), .B(n1808), .ZN(N4586) );
  aoi22d1 U2721 ( .A1(n1818), .A2(spi_master_mosi[2]), .B1(n1821), .B2(
        csrbank9_control0_w[2]), .ZN(n1811) );
  aoi22d1 U2722 ( .A1(n4579), .A2(csrbank9_cs0_w[2]), .B1(n1822), .B2(
        spi_master_miso_status[2]), .ZN(n1810) );
  oai211d1 U2723 ( .C1(n1827), .C2(n3065), .A(n1811), .B(n1810), .ZN(N4587) );
  aoi22d1 U2724 ( .A1(n1818), .A2(spi_master_mosi[3]), .B1(n1821), .B2(
        csrbank9_control0_w[3]), .ZN(n1813) );
  aoi22d1 U2725 ( .A1(n4579), .A2(csrbank9_cs0_w[3]), .B1(n1822), .B2(
        spi_master_miso_status[3]), .ZN(n1812) );
  oai211d1 U2726 ( .C1(n1827), .C2(n3066), .A(n1813), .B(n1812), .ZN(N4588) );
  aoi22d1 U2727 ( .A1(n4579), .A2(csrbank9_cs0_w[4]), .B1(n1822), .B2(
        spi_master_miso_status[4]), .ZN(n1815) );
  aoi22d1 U2728 ( .A1(n1818), .A2(spi_master_mosi[4]), .B1(n1821), .B2(
        csrbank9_control0_w[4]), .ZN(n1814) );
  oai211d1 U2729 ( .C1(n1827), .C2(n3067), .A(n1815), .B(n1814), .ZN(N4589) );
  aoi22d1 U2730 ( .A1(n1821), .A2(csrbank9_control0_w[5]), .B1(n1822), .B2(
        spi_master_miso_status[5]), .ZN(n1817) );
  aoi22d1 U2731 ( .A1(n1818), .A2(spi_master_mosi[5]), .B1(n4579), .B2(
        csrbank9_cs0_w[5]), .ZN(n1816) );
  oai211d1 U2732 ( .C1(n1827), .C2(n3068), .A(n1817), .B(n1816), .ZN(N4590) );
  inv0d0 U2733 ( .I(n1818), .ZN(n1825) );
  inv0d0 U2734 ( .I(spi_master_mosi[6]), .ZN(n4563) );
  inv0d0 U2735 ( .I(n1827), .ZN(n3063) );
  aoi22d1 U2736 ( .A1(n3063), .A2(spi_master_clk_divider0[6]), .B1(n1822), 
        .B2(spi_master_miso_status[6]), .ZN(n1820) );
  aoi22d1 U2737 ( .A1(n1821), .A2(csrbank9_control0_w[6]), .B1(n4579), .B2(
        csrbank9_cs0_w[6]), .ZN(n1819) );
  oai211d1 U2738 ( .C1(n1825), .C2(n4563), .A(n1820), .B(n1819), .ZN(N4591) );
  inv0d0 U2739 ( .I(spi_master_mosi[7]), .ZN(n4567) );
  aoi22d1 U2740 ( .A1(n3063), .A2(spi_master_clk_divider0[7]), .B1(n1821), 
        .B2(csrbank9_control0_w[7]), .ZN(n1824) );
  aoi22d1 U2741 ( .A1(n4579), .A2(csrbank9_cs0_w[7]), .B1(n1822), .B2(
        spi_master_miso_status[7]), .ZN(n1823) );
  oai211d1 U2742 ( .C1(n1825), .C2(n4567), .A(n1824), .B(n1823), .ZN(N4592) );
  inv0d0 U2743 ( .I(csrbank9_cs0_w[8]), .ZN(n4591) );
  inv0d0 U2744 ( .I(spi_master_length0[0]), .ZN(n4635) );
  oai222d1 U2745 ( .A1(n4591), .A2(n1828), .B1(n3072), .B2(n1827), .C1(n1826), 
        .C2(n4635), .ZN(N4593) );
  inv0d0 U2746 ( .I(csrbank9_cs0_w[9]), .ZN(n4592) );
  inv0d0 U2747 ( .I(spi_master_length0[1]), .ZN(n4636) );
  oai222d1 U2748 ( .A1(n4592), .A2(n1828), .B1(n3073), .B2(n1827), .C1(n1826), 
        .C2(n4636), .ZN(N4594) );
  inv0d0 U2749 ( .I(csrbank9_cs0_w[10]), .ZN(n4594) );
  inv0d0 U2750 ( .I(spi_master_length0[2]), .ZN(n4637) );
  oai222d1 U2751 ( .A1(n4594), .A2(n1828), .B1(n3074), .B2(n1827), .C1(n1826), 
        .C2(n4637), .ZN(N4595) );
  inv0d0 U2752 ( .I(csrbank9_cs0_w[11]), .ZN(n4596) );
  inv0d0 U2753 ( .I(spi_master_length0[3]), .ZN(n4638) );
  oai222d1 U2754 ( .A1(n4596), .A2(n1828), .B1(n3075), .B2(n1827), .C1(n1826), 
        .C2(n4638), .ZN(N4596) );
  inv0d0 U2755 ( .I(csrbank9_cs0_w[12]), .ZN(n4597) );
  inv0d0 U2756 ( .I(spi_master_length0[4]), .ZN(n4639) );
  oai222d1 U2757 ( .A1(n4597), .A2(n1828), .B1(n3076), .B2(n1827), .C1(n1826), 
        .C2(n4639), .ZN(N4597) );
  inv0d0 U2758 ( .I(csrbank9_cs0_w[13]), .ZN(n4599) );
  inv0d0 U2759 ( .I(spi_master_length0[5]), .ZN(n4640) );
  oai222d1 U2760 ( .A1(n4599), .A2(n1828), .B1(n3077), .B2(n1827), .C1(n1826), 
        .C2(n4640), .ZN(N4598) );
  inv0d0 U2761 ( .I(csrbank9_cs0_w[14]), .ZN(n4600) );
  inv0d0 U2762 ( .I(spi_master_length0[6]), .ZN(n4641) );
  oai222d1 U2763 ( .A1(n4600), .A2(n1828), .B1(n3078), .B2(n1827), .C1(n1826), 
        .C2(n4641), .ZN(N4599) );
  inv0d0 U2764 ( .I(csrbank9_cs0_w[15]), .ZN(n4602) );
  inv0d0 U2765 ( .I(spi_master_length0[7]), .ZN(n4642) );
  oai222d1 U2766 ( .A1(n4602), .A2(n1828), .B1(n3079), .B2(n1827), .C1(n1826), 
        .C2(n4642), .ZN(N4600) );
  aoi22d1 U2767 ( .A1(n4998), .A2(gpio_mode1_pad), .B1(n1839), .B2(
        csrbank5_in_w), .ZN(n1833) );
  aoi22d1 U2768 ( .A1(n1902), .A2(n6130), .B1(n4952), .B2(csrbank5_ien0_w), 
        .ZN(n1832) );
  aoi22d1 U2769 ( .A1(n1838), .A2(csrbank5_oe0_w), .B1(n2457), .B2(
        gpio_mode0_pad), .ZN(n1831) );
  inv0d0 U2770 ( .I(n1829), .ZN(n3058) );
  nr02d0 U2771 ( .A1(n3058), .A2(n2469), .ZN(n2450) );
  nd02d0 U2772 ( .A1(n1903), .A2(n2450), .ZN(n1830) );
  aoi31d1 U2773 ( .B1(n1833), .B2(n1832), .B3(n1831), .A(n1830), .ZN(N4331) );
  inv0d0 U2774 ( .I(csrbank5_ien0_w), .ZN(gpio_inenb_pad) );
  oai21d1 U2775 ( .B1(n4685), .B2(n1834), .A(
        mgmtsoc_port_master_user_port_sink_valid), .ZN(n4724) );
  aoi22d1 U2776 ( .A1(n4998), .A2(mgmtsoc_litespimmap_spi_dummy_bits[0]), .B1(
        n1839), .B2(n4724), .ZN(n1837) );
  inv0d0 U2777 ( .I(mgmtsoc_master_rxtx_w[0]), .ZN(n4687) );
  inv0d0 U2778 ( .I(mgmtsoc_master_tx_fifo_sink_payload_len[0]), .ZN(n4774) );
  oai22d1 U2779 ( .A1(n2451), .A2(n4687), .B1(n2454), .B2(n4774), .ZN(n1835)
         );
  aoi21d1 U2780 ( .B1(n2457), .B2(\litespi_request[1] ), .A(n1835), .ZN(n1836)
         );
  aoi21d1 U2781 ( .B1(n1837), .B2(n1836), .A(n1840), .ZN(N4243) );
  aoi22d1 U2782 ( .A1(n1838), .A2(mgmtsoc_master_rxtx_w[1]), .B1(n4952), .B2(
        mgmtsoc_master_tx_fifo_sink_payload_len[1]), .ZN(n1842) );
  aoi22d1 U2783 ( .A1(n4998), .A2(mgmtsoc_litespimmap_spi_dummy_bits[1]), .B1(
        \mgmtsoc_master_status_status[1] ), .B2(n1839), .ZN(n1841) );
  aoi21d1 U2784 ( .B1(n1842), .B2(n1841), .A(n1840), .ZN(N4244) );
  inv0d0 U2785 ( .I(mgmtsoc_master_tx_fifo_sink_payload_len[2]), .ZN(n4776) );
  buffd1 U2786 ( .I(n1844), .Z(n4773) );
  inv0d0 U2787 ( .I(mgmtsoc_master_rxtx_w[2]), .ZN(n4689) );
  inv0d0 U2788 ( .I(mgmtsoc_litespimmap_spi_dummy_bits[2]), .ZN(n4814) );
  oai222d1 U2789 ( .A1(n4776), .A2(n4773), .B1(n4689), .B2(n1845), .C1(n4814), 
        .C2(n4810), .ZN(N4245) );
  inv0d0 U2790 ( .I(mgmtsoc_master_tx_fifo_sink_payload_len[3]), .ZN(n4777) );
  inv0d0 U2791 ( .I(mgmtsoc_master_rxtx_w[3]), .ZN(n4690) );
  oai222d1 U2792 ( .A1(n4777), .A2(n1844), .B1(n4690), .B2(n4723), .C1(n4815), 
        .C2(n4810), .ZN(N4246) );
  inv0d0 U2793 ( .I(mgmtsoc_master_tx_fifo_sink_payload_len[4]), .ZN(n4778) );
  inv0d0 U2794 ( .I(mgmtsoc_master_rxtx_w[4]), .ZN(n4691) );
  oai222d1 U2795 ( .A1(n4778), .A2(n1844), .B1(n4691), .B2(n1845), .C1(n4816), 
        .C2(n4810), .ZN(N4247) );
  inv0d0 U2796 ( .I(mgmtsoc_master_tx_fifo_sink_payload_len[5]), .ZN(n4779) );
  inv0d0 U2797 ( .I(mgmtsoc_master_rxtx_w[5]), .ZN(n4692) );
  oai222d1 U2798 ( .A1(n4779), .A2(n1844), .B1(n4692), .B2(n4723), .C1(n4817), 
        .C2(n4810), .ZN(N4248) );
  inv0d0 U2799 ( .I(mgmtsoc_master_len[6]), .ZN(n4780) );
  inv0d0 U2800 ( .I(mgmtsoc_master_rxtx_w[6]), .ZN(n4693) );
  oai222d1 U2801 ( .A1(n4780), .A2(n1844), .B1(n4693), .B2(n4723), .C1(n4810), 
        .C2(n4818), .ZN(N4249) );
  inv0d0 U2802 ( .I(mgmtsoc_master_len[7]), .ZN(n4781) );
  inv0d0 U2803 ( .I(mgmtsoc_master_rxtx_w[7]), .ZN(n4694) );
  inv0d0 U2804 ( .I(mgmtsoc_litespimmap_spi_dummy_bits[7]), .ZN(n4820) );
  oai222d1 U2805 ( .A1(n4781), .A2(n4773), .B1(n4694), .B2(n4723), .C1(n4810), 
        .C2(n4820), .ZN(N4250) );
  inv0d0 U2806 ( .I(mgmtsoc_master_rxtx_w[8]), .ZN(n4695) );
  inv0d0 U2807 ( .I(mgmtsoc_master_tx_fifo_sink_payload_width[0]), .ZN(n4782)
         );
  oai22d1 U2808 ( .A1(n4723), .A2(n4695), .B1(n4773), .B2(n4782), .ZN(N4251)
         );
  inv0d0 U2809 ( .I(mgmtsoc_master_rxtx_w[9]), .ZN(n4696) );
  inv0d0 U2810 ( .I(mgmtsoc_master_tx_fifo_sink_payload_width[1]), .ZN(n4784)
         );
  oai22d1 U2811 ( .A1(n1845), .A2(n4696), .B1(n4773), .B2(n4784), .ZN(N4252)
         );
  inv0d0 U2812 ( .I(mgmtsoc_master_rxtx_w[10]), .ZN(n4697) );
  inv0d0 U2813 ( .I(mgmtsoc_master_tx_fifo_sink_payload_width[2]), .ZN(n4785)
         );
  oai22d1 U2814 ( .A1(n4723), .A2(n4697), .B1(n1844), .B2(n4785), .ZN(N4253)
         );
  inv0d0 U2815 ( .I(mgmtsoc_master_rxtx_w[11]), .ZN(n4698) );
  inv0d0 U2816 ( .I(mgmtsoc_master_tx_fifo_sink_payload_width[3]), .ZN(n4786)
         );
  oai22d1 U2817 ( .A1(n4723), .A2(n4698), .B1(n4773), .B2(n4786), .ZN(N4254)
         );
  inv0d0 U2818 ( .I(mgmtsoc_master_rxtx_w[12]), .ZN(n4699) );
  inv0d0 U2819 ( .I(csrbank3_master_phyconfig0_w[12]), .ZN(n4788) );
  oai22d1 U2820 ( .A1(n4723), .A2(n4699), .B1(n1844), .B2(n4788), .ZN(N4255)
         );
  inv0d0 U2821 ( .I(mgmtsoc_master_rxtx_w[13]), .ZN(n4700) );
  inv0d0 U2822 ( .I(csrbank3_master_phyconfig0_w[13]), .ZN(n4789) );
  oai22d1 U2823 ( .A1(n4723), .A2(n4700), .B1(n1844), .B2(n4789), .ZN(N4256)
         );
  inv0d0 U2824 ( .I(mgmtsoc_master_rxtx_w[14]), .ZN(n4701) );
  inv0d0 U2825 ( .I(csrbank3_master_phyconfig0_w[14]), .ZN(n4791) );
  oai22d1 U2826 ( .A1(n1845), .A2(n4701), .B1(n4773), .B2(n4791), .ZN(N4257)
         );
  inv0d0 U2827 ( .I(mgmtsoc_master_rxtx_w[15]), .ZN(n4702) );
  inv0d0 U2828 ( .I(csrbank3_master_phyconfig0_w[15]), .ZN(n4792) );
  oai22d1 U2829 ( .A1(n1845), .A2(n4702), .B1(n1844), .B2(n4792), .ZN(N4258)
         );
  inv0d0 U2830 ( .I(mgmtsoc_master_rxtx_w[16]), .ZN(n4703) );
  inv0d0 U2831 ( .I(mgmtsoc_master_tx_fifo_sink_payload_mask[0]), .ZN(n4794)
         );
  oai22d1 U2832 ( .A1(n1845), .A2(n4703), .B1(n4773), .B2(n4794), .ZN(N4259)
         );
  inv0d0 U2833 ( .I(mgmtsoc_master_rxtx_w[17]), .ZN(n4704) );
  inv0d0 U2834 ( .I(mgmtsoc_master_tx_fifo_sink_payload_mask[1]), .ZN(n4796)
         );
  oai22d1 U2835 ( .A1(n1845), .A2(n4704), .B1(n4773), .B2(n4796), .ZN(N4260)
         );
  inv0d0 U2836 ( .I(mgmtsoc_master_rxtx_w[18]), .ZN(n4705) );
  inv0d0 U2837 ( .I(mgmtsoc_master_tx_fifo_sink_payload_mask[2]), .ZN(n4798)
         );
  oai22d1 U2838 ( .A1(n4723), .A2(n4705), .B1(n4773), .B2(n4798), .ZN(N4261)
         );
  inv0d0 U2839 ( .I(mgmtsoc_master_rxtx_w[19]), .ZN(n4706) );
  inv0d0 U2840 ( .I(mgmtsoc_master_tx_fifo_sink_payload_mask[3]), .ZN(n4799)
         );
  oai22d1 U2841 ( .A1(n4723), .A2(n4706), .B1(n4773), .B2(n4799), .ZN(N4262)
         );
  inv0d0 U2842 ( .I(mgmtsoc_master_rxtx_w[20]), .ZN(n4707) );
  inv0d0 U2843 ( .I(mgmtsoc_master_tx_fifo_sink_payload_mask[4]), .ZN(n4800)
         );
  oai22d1 U2844 ( .A1(n4723), .A2(n4707), .B1(n4773), .B2(n4800), .ZN(N4263)
         );
  inv0d0 U2845 ( .I(mgmtsoc_master_rxtx_w[21]), .ZN(n4708) );
  inv0d0 U2846 ( .I(mgmtsoc_master_tx_fifo_sink_payload_mask[5]), .ZN(n4801)
         );
  oai22d1 U2847 ( .A1(n4723), .A2(n4708), .B1(n4773), .B2(n4801), .ZN(N4264)
         );
  inv0d0 U2848 ( .I(mgmtsoc_master_rxtx_w[22]), .ZN(n4709) );
  inv0d0 U2849 ( .I(mgmtsoc_master_tx_fifo_sink_payload_mask[6]), .ZN(n4802)
         );
  oai22d1 U2850 ( .A1(n4723), .A2(n4709), .B1(n4773), .B2(n4802), .ZN(N4265)
         );
  inv0d0 U2851 ( .I(mgmtsoc_master_rxtx_w[23]), .ZN(n4710) );
  inv0d0 U2852 ( .I(mgmtsoc_master_tx_fifo_sink_payload_mask[7]), .ZN(n4803)
         );
  oai22d1 U2853 ( .A1(n4723), .A2(n4710), .B1(n4773), .B2(n4803), .ZN(N4266)
         );
  nd12d1 U2854 ( .A1(n1846), .A2(n5241), .ZN(n1860) );
  buffd1 U2855 ( .I(n1860), .Z(n1865) );
  inv0d0 U2856 ( .I(mgmtsoc_bus_errors_status[0]), .ZN(n5113) );
  inv0d0 U2857 ( .I(csrbank0_reset0_w[0]), .ZN(n5289) );
  inv0d0 U2858 ( .I(csrbank0_scratch0_w[0]), .ZN(n5242) );
  nd12d1 U2859 ( .A1(n1847), .A2(n5241), .ZN(n1863) );
  buffd1 U2860 ( .I(n1863), .Z(n1864) );
  oai222d1 U2861 ( .A1(n1865), .A2(n5113), .B1(n5289), .B2(n1848), .C1(n5242), 
        .C2(n1864), .ZN(N4099) );
  inv0d0 U2862 ( .I(csrbank0_scratch0_w[1]), .ZN(n5243) );
  inv0d0 U2863 ( .I(csrbank0_reset0_w[1]), .ZN(n5292) );
  inv0d0 U2864 ( .I(mgmtsoc_bus_errors_status[1]), .ZN(n5239) );
  oai222d1 U2865 ( .A1(n5243), .A2(n1864), .B1(n5292), .B2(n1848), .C1(n5239), 
        .C2(n1860), .ZN(N4100) );
  inv0d0 U2866 ( .I(mgmtsoc_bus_errors_status[2]), .ZN(n5234) );
  inv0d0 U2867 ( .I(csrbank0_scratch0_w[2]), .ZN(n5244) );
  oai22d1 U2868 ( .A1(n1860), .A2(n5234), .B1(n1864), .B2(n5244), .ZN(N4101)
         );
  inv0d0 U2869 ( .I(mgmtsoc_bus_errors_status[3]), .ZN(n5230) );
  inv0d0 U2870 ( .I(csrbank0_scratch0_w[3]), .ZN(n1849) );
  oai22d1 U2871 ( .A1(n1860), .A2(n5230), .B1(n1864), .B2(n1849), .ZN(N4102)
         );
  inv0d0 U2872 ( .I(mgmtsoc_bus_errors_status[4]), .ZN(n5226) );
  inv0d0 U2873 ( .I(csrbank0_scratch0_w[4]), .ZN(n1850) );
  oai22d1 U2874 ( .A1(n1860), .A2(n5226), .B1(n1864), .B2(n1850), .ZN(N4103)
         );
  inv0d0 U2875 ( .I(mgmtsoc_bus_errors_status[5]), .ZN(n5222) );
  inv0d0 U2876 ( .I(csrbank0_scratch0_w[5]), .ZN(n1851) );
  oai22d1 U2877 ( .A1(n1865), .A2(n5222), .B1(n1863), .B2(n1851), .ZN(N4104)
         );
  inv0d0 U2878 ( .I(mgmtsoc_bus_errors_status[6]), .ZN(n5218) );
  inv0d0 U2879 ( .I(csrbank0_scratch0_w[6]), .ZN(n1852) );
  oai22d1 U2880 ( .A1(n1860), .A2(n5218), .B1(n1863), .B2(n1852), .ZN(N4105)
         );
  inv0d0 U2881 ( .I(mgmtsoc_bus_errors_status[7]), .ZN(n5213) );
  inv0d0 U2882 ( .I(csrbank0_scratch0_w[7]), .ZN(n5250) );
  oai22d1 U2883 ( .A1(n1860), .A2(n5213), .B1(n1863), .B2(n5250), .ZN(N4106)
         );
  inv0d0 U2884 ( .I(mgmtsoc_bus_errors_status[8]), .ZN(n5209) );
  inv0d0 U2885 ( .I(csrbank0_scratch0_w[8]), .ZN(n5252) );
  oai22d1 U2886 ( .A1(n1860), .A2(n5209), .B1(n1863), .B2(n5252), .ZN(N4107)
         );
  inv0d0 U2887 ( .I(mgmtsoc_bus_errors_status[9]), .ZN(n5205) );
  inv0d0 U2888 ( .I(csrbank0_scratch0_w[9]), .ZN(n1853) );
  oai22d1 U2889 ( .A1(n1860), .A2(n5205), .B1(n1864), .B2(n1853), .ZN(N4108)
         );
  inv0d0 U2890 ( .I(mgmtsoc_bus_errors_status[10]), .ZN(n5200) );
  inv0d0 U2891 ( .I(csrbank0_scratch0_w[10]), .ZN(n1854) );
  oai22d1 U2892 ( .A1(n1865), .A2(n5200), .B1(n1863), .B2(n1854), .ZN(N4109)
         );
  inv0d0 U2893 ( .I(mgmtsoc_bus_errors_status[11]), .ZN(n5196) );
  inv0d0 U2894 ( .I(csrbank0_scratch0_w[11]), .ZN(n5253) );
  oai22d1 U2895 ( .A1(n1860), .A2(n5196), .B1(n1864), .B2(n5253), .ZN(N4110)
         );
  inv0d0 U2896 ( .I(mgmtsoc_bus_errors_status[12]), .ZN(n5192) );
  inv0d0 U2897 ( .I(csrbank0_scratch0_w[12]), .ZN(n1855) );
  oai22d1 U2898 ( .A1(n1860), .A2(n5192), .B1(n1863), .B2(n1855), .ZN(N4111)
         );
  inv0d0 U2899 ( .I(mgmtsoc_bus_errors_status[13]), .ZN(n5188) );
  inv0d0 U2900 ( .I(csrbank0_scratch0_w[13]), .ZN(n5255) );
  oai22d1 U2901 ( .A1(n1860), .A2(n5188), .B1(n1863), .B2(n5255), .ZN(N4112)
         );
  inv0d0 U2902 ( .I(mgmtsoc_bus_errors_status[14]), .ZN(n5184) );
  inv0d0 U2903 ( .I(csrbank0_scratch0_w[14]), .ZN(n1856) );
  oai22d1 U2904 ( .A1(n1860), .A2(n5184), .B1(n1863), .B2(n1856), .ZN(N4113)
         );
  inv0d0 U2905 ( .I(mgmtsoc_bus_errors_status[15]), .ZN(n5180) );
  inv0d0 U2906 ( .I(csrbank0_scratch0_w[15]), .ZN(n5256) );
  oai22d1 U2907 ( .A1(n1860), .A2(n5180), .B1(n1863), .B2(n5256), .ZN(N4114)
         );
  inv0d0 U2908 ( .I(mgmtsoc_bus_errors_status[16]), .ZN(n5176) );
  inv0d0 U2909 ( .I(csrbank0_scratch0_w[16]), .ZN(n5257) );
  oai22d1 U2910 ( .A1(n1865), .A2(n5176), .B1(n1863), .B2(n5257), .ZN(N4115)
         );
  inv0d0 U2911 ( .I(mgmtsoc_bus_errors_status[17]), .ZN(n5172) );
  inv0d0 U2912 ( .I(csrbank0_scratch0_w[17]), .ZN(n5258) );
  oai22d1 U2913 ( .A1(n1865), .A2(n5172), .B1(n1864), .B2(n5258), .ZN(N4116)
         );
  inv0d0 U2914 ( .I(mgmtsoc_bus_errors_status[18]), .ZN(n5168) );
  inv0d0 U2915 ( .I(csrbank0_scratch0_w[18]), .ZN(n1857) );
  oai22d1 U2916 ( .A1(n1865), .A2(n5168), .B1(n1863), .B2(n1857), .ZN(N4117)
         );
  inv0d0 U2917 ( .I(mgmtsoc_bus_errors_status[19]), .ZN(n5164) );
  inv0d0 U2918 ( .I(csrbank0_scratch0_w[19]), .ZN(n5261) );
  oai22d1 U2919 ( .A1(n1860), .A2(n5164), .B1(n1864), .B2(n5261), .ZN(N4118)
         );
  inv0d0 U2920 ( .I(mgmtsoc_bus_errors_status[20]), .ZN(n5160) );
  inv0d0 U2921 ( .I(csrbank0_scratch0_w[20]), .ZN(n1858) );
  oai22d1 U2922 ( .A1(n1865), .A2(n5160), .B1(n1863), .B2(n1858), .ZN(N4119)
         );
  inv0d0 U2923 ( .I(mgmtsoc_bus_errors_status[21]), .ZN(n5156) );
  inv0d0 U2924 ( .I(csrbank0_scratch0_w[21]), .ZN(n1859) );
  oai22d1 U2925 ( .A1(n1865), .A2(n5156), .B1(n1864), .B2(n1859), .ZN(N4120)
         );
  inv0d0 U2926 ( .I(mgmtsoc_bus_errors_status[22]), .ZN(n5152) );
  inv0d0 U2927 ( .I(csrbank0_scratch0_w[22]), .ZN(n5265) );
  oai22d1 U2928 ( .A1(n1860), .A2(n5152), .B1(n1864), .B2(n5265), .ZN(N4121)
         );
  inv0d0 U2929 ( .I(mgmtsoc_bus_errors_status[23]), .ZN(n5148) );
  inv0d0 U2930 ( .I(csrbank0_scratch0_w[23]), .ZN(n5267) );
  oai22d1 U2931 ( .A1(n1865), .A2(n5148), .B1(n1864), .B2(n5267), .ZN(N4122)
         );
  inv0d0 U2932 ( .I(mgmtsoc_bus_errors_status[24]), .ZN(n5144) );
  inv0d0 U2933 ( .I(csrbank0_scratch0_w[24]), .ZN(n5269) );
  oai22d1 U2934 ( .A1(n1865), .A2(n5144), .B1(n1863), .B2(n5269), .ZN(N4123)
         );
  inv0d0 U2935 ( .I(mgmtsoc_bus_errors_status[25]), .ZN(n5140) );
  inv0d0 U2936 ( .I(csrbank0_scratch0_w[25]), .ZN(n1861) );
  oai22d1 U2937 ( .A1(n1865), .A2(n5140), .B1(n1863), .B2(n1861), .ZN(N4124)
         );
  inv0d0 U2938 ( .I(mgmtsoc_bus_errors_status[26]), .ZN(n5136) );
  inv0d0 U2939 ( .I(csrbank0_scratch0_w[26]), .ZN(n5272) );
  oai22d1 U2940 ( .A1(n1865), .A2(n5136), .B1(n1864), .B2(n5272), .ZN(N4125)
         );
  inv0d0 U2941 ( .I(mgmtsoc_bus_errors_status[27]), .ZN(n5132) );
  inv0d0 U2942 ( .I(csrbank0_scratch0_w[27]), .ZN(n5274) );
  oai22d1 U2943 ( .A1(n1865), .A2(n5132), .B1(n1864), .B2(n5274), .ZN(N4126)
         );
  inv0d0 U2944 ( .I(mgmtsoc_bus_errors_status[28]), .ZN(n5128) );
  inv0d0 U2945 ( .I(csrbank0_scratch0_w[28]), .ZN(n1862) );
  oai22d1 U2946 ( .A1(n1865), .A2(n5128), .B1(n1863), .B2(n1862), .ZN(N4127)
         );
  inv0d0 U2947 ( .I(mgmtsoc_bus_errors_status[29]), .ZN(n5124) );
  inv0d0 U2948 ( .I(csrbank0_scratch0_w[29]), .ZN(n5278) );
  oai22d1 U2949 ( .A1(n1865), .A2(n5124), .B1(n1864), .B2(n5278), .ZN(N4128)
         );
  inv0d0 U2950 ( .I(mgmtsoc_bus_errors_status[30]), .ZN(n5120) );
  inv0d0 U2951 ( .I(csrbank0_scratch0_w[30]), .ZN(n5281) );
  oai22d1 U2952 ( .A1(n1865), .A2(n5120), .B1(n1864), .B2(n5281), .ZN(N4129)
         );
  inv0d0 U2953 ( .I(mgmtsoc_bus_errors_status[31]), .ZN(n5116) );
  inv0d0 U2954 ( .I(csrbank0_scratch0_w[31]), .ZN(n5284) );
  oai22d1 U2955 ( .A1(n1865), .A2(n5116), .B1(n1864), .B2(n5284), .ZN(N4130)
         );
  inv0d0 U2956 ( .I(mgmtsoc_litespisdrphycore_sr_out[28]), .ZN(n5815) );
  inv0d0 U2957 ( .I(mgmtsoc_litespisdrphycore_sr_out[30]), .ZN(n5799) );
  inv0d0 U2958 ( .I(mgmtsoc_litespisdrphycore_sr_out[24]), .ZN(n5859) );
  oai22d1 U2959 ( .A1(n1867), .A2(n5799), .B1(n1866), .B2(n5859), .ZN(n1868)
         );
  aoi21d1 U2960 ( .B1(mgmtsoc_litespisdrphycore_sr_out[31]), .B2(n5736), .A(
        n1868), .ZN(n1869) );
  oai21d1 U2961 ( .B1(n1870), .B2(n5815), .A(n1869), .ZN(
        mgmtsoc_litespisdrphycore_dq_o) );
  aoi22d1 U2962 ( .A1(litespi_tx_mux_sel), .A2(
        \mgmtsoc_port_master_user_port_sink_payload_mask[0] ), .B1(n1871), 
        .B2(n4840), .ZN(n4547) );
  inv0d0 U2963 ( .I(uart_rx_fifo_rdport_adr[3]), .ZN(n1873) );
  inv0d0 U2964 ( .I(uart_rx_fifo_rdport_adr[1]), .ZN(n2511) );
  nr03d0 U2965 ( .A1(uart_rx_fifo_rdport_adr[2]), .A2(n1873), .A3(n2511), .ZN(
        n2984) );
  nr03d0 U2966 ( .A1(uart_rx_fifo_rdport_adr[3]), .A2(
        uart_rx_fifo_rdport_adr[2]), .A3(n2511), .ZN(n2959) );
  aoi22d1 U2967 ( .A1(\storage_1[11][0] ), .A2(n2984), .B1(\storage_1[3][0] ), 
        .B2(n2959), .ZN(n1884) );
  inv0d0 U2968 ( .I(\storage_1[15][0] ), .ZN(n2891) );
  nd02d0 U2969 ( .A1(uart_rx_fifo_rdport_adr[1]), .A2(
        uart_rx_fifo_rdport_adr[2]), .ZN(n2512) );
  nr02d1 U2970 ( .A1(n1873), .A2(n2512), .ZN(n3033) );
  inv0d0 U2971 ( .I(n3033), .ZN(n3003) );
  inv0d0 U2972 ( .I(\storage_1[9][0] ), .ZN(n2904) );
  nr03d0 U2973 ( .A1(uart_rx_fifo_rdport_adr[1]), .A2(
        uart_rx_fifo_rdport_adr[2]), .A3(n1873), .ZN(n3013) );
  buffd1 U2974 ( .I(n3013), .Z(n3034) );
  inv0d0 U2975 ( .I(n3034), .ZN(n3001) );
  oai22d1 U2976 ( .A1(n2891), .A2(n3003), .B1(n2904), .B2(n3001), .ZN(n1876)
         );
  inv0d0 U2977 ( .I(\storage_1[5][0] ), .ZN(n2918) );
  inv0d0 U2978 ( .I(uart_rx_fifo_rdport_adr[2]), .ZN(n1872) );
  nr03d0 U2979 ( .A1(uart_rx_fifo_rdport_adr[1]), .A2(
        uart_rx_fifo_rdport_adr[3]), .A3(n1872), .ZN(n3031) );
  buffd1 U2980 ( .I(n3031), .Z(n3012) );
  inv0d0 U2981 ( .I(n3012), .ZN(n2999) );
  inv0d0 U2982 ( .I(\storage_1[1][0] ), .ZN(n2927) );
  nr03d0 U2983 ( .A1(uart_rx_fifo_rdport_adr[1]), .A2(
        uart_rx_fifo_rdport_adr[3]), .A3(uart_rx_fifo_rdport_adr[2]), .ZN(
        n2958) );
  buffd1 U2984 ( .I(n2958), .Z(n3030) );
  inv0d0 U2985 ( .I(n3030), .ZN(n2997) );
  oai22d1 U2986 ( .A1(n2918), .A2(n2999), .B1(n2927), .B2(n2997), .ZN(n1875)
         );
  inv0d0 U2987 ( .I(\storage_1[13][0] ), .ZN(n2895) );
  nr03d0 U2988 ( .A1(uart_rx_fifo_rdport_adr[1]), .A2(n1873), .A3(n1872), .ZN(
        n2985) );
  buffd1 U2989 ( .I(n2985), .Z(n3037) );
  inv0d0 U2990 ( .I(n3037), .ZN(n3007) );
  inv0d0 U2991 ( .I(\storage_1[7][0] ), .ZN(n2910) );
  nr02d1 U2992 ( .A1(uart_rx_fifo_rdport_adr[3]), .A2(n2512), .ZN(n3036) );
  inv0d0 U2993 ( .I(n3036), .ZN(n3005) );
  oai22d1 U2994 ( .A1(n2895), .A2(n3007), .B1(n2910), .B2(n3005), .ZN(n1874)
         );
  nr03d0 U2995 ( .A1(n1876), .A2(n1875), .A3(n1874), .ZN(n1883) );
  inv0d0 U2996 ( .I(uart_rx_fifo_level0[4]), .ZN(n2549) );
  nd02d0 U2997 ( .A1(uart_pending_r[1]), .A2(uart_pending_re), .ZN(n2660) );
  nd02d0 U2998 ( .A1(\uart_status_status[1] ), .A2(n2660), .ZN(n2548) );
  oaim21d1 U2999 ( .B1(n2549), .B2(n2550), .A(n2548), .ZN(n3020) );
  inv0d1 U3000 ( .I(n3020), .ZN(n3046) );
  nd02d0 U3001 ( .A1(n3046), .A2(uart_rx_fifo_rdport_adr[0]), .ZN(n3022) );
  nr02d0 U3002 ( .A1(uart_rx_fifo_rdport_adr[0]), .A2(n3020), .ZN(n3019) );
  aoi22d1 U3003 ( .A1(\storage_1[8][0] ), .A2(n3013), .B1(\storage_1[6][0] ), 
        .B2(n3036), .ZN(n1880) );
  aoi22d1 U3004 ( .A1(\storage_1[14][0] ), .A2(n3033), .B1(\storage_1[4][0] ), 
        .B2(n3031), .ZN(n1879) );
  buffd1 U3005 ( .I(n2959), .Z(n3032) );
  aoi22d1 U3006 ( .A1(\storage_1[2][0] ), .A2(n3032), .B1(\storage_1[0][0] ), 
        .B2(n2958), .ZN(n1878) );
  buffd1 U3007 ( .I(n2984), .Z(n3035) );
  aoi22d1 U3008 ( .A1(\storage_1[12][0] ), .A2(n2985), .B1(\storage_1[10][0] ), 
        .B2(n3035), .ZN(n1877) );
  aoi22d1 U3009 ( .A1(uart_rx_fifo_fifo_out_payload_data[0]), .A2(n3020), .B1(
        n3019), .B2(n1881), .ZN(n1882) );
  aon211d1 U3010 ( .C1(n1884), .C2(n1883), .B(n3022), .A(n1882), .ZN(n4546) );
  an02d0 U3011 ( .A1(n2013), .A2(mprj_dat_o[0]), .Z(n4582) );
  inv0d2 U3012 ( .I(n4582), .ZN(n5290) );
  inv0d0 U3013 ( .I(spi_master_mosi[0]), .ZN(n4553) );
  inv0d0 U3014 ( .I(n1886), .ZN(n1885) );
  aoi22d1 U3015 ( .A1(n1886), .A2(n5290), .B1(n4553), .B2(n1885), .ZN(n4545)
         );
  nd02d0 U3016 ( .A1(n2013), .A2(mprj_dat_o[1]), .ZN(n2639) );
  buffd1 U3017 ( .I(n2639), .Z(n4862) );
  buffd1 U3018 ( .I(n4862), .Z(n5294) );
  inv0d0 U3019 ( .I(spi_master_mosi[1]), .ZN(n4555) );
  aoi22d1 U3020 ( .A1(n1886), .A2(n5294), .B1(n4555), .B2(n1885), .ZN(n4544)
         );
  nd02d0 U3021 ( .A1(n2013), .A2(mprj_dat_o[2]), .ZN(n5245) );
  buffd3 U3022 ( .I(n5245), .Z(n5004) );
  inv0d0 U3023 ( .I(spi_master_mosi[2]), .ZN(n4556) );
  aoi22d1 U3024 ( .A1(n1886), .A2(n5004), .B1(n4556), .B2(n1885), .ZN(n4543)
         );
  inv0d0 U3025 ( .I(spi_master_mosi[3]), .ZN(n4557) );
  aoi22d1 U3026 ( .A1(n1886), .A2(n2625), .B1(n4557), .B2(n1885), .ZN(n4542)
         );
  buffd1 U3027 ( .I(n4866), .Z(n5008) );
  inv0d0 U3028 ( .I(spi_master_mosi[4]), .ZN(n4559) );
  aoi22d1 U3029 ( .A1(n1886), .A2(n5008), .B1(n4559), .B2(n1885), .ZN(n4541)
         );
  buffd1 U3030 ( .I(n2640), .Z(n5010) );
  inv0d0 U3031 ( .I(spi_master_mosi[5]), .ZN(n4561) );
  aoi22d1 U3032 ( .A1(n1886), .A2(n5010), .B1(n4561), .B2(n1885), .ZN(n4540)
         );
  nd02d0 U3033 ( .A1(n2013), .A2(mprj_dat_o[6]), .ZN(n2641) );
  buffd1 U3034 ( .I(n2641), .Z(n5012) );
  aoi22d1 U3035 ( .A1(n1886), .A2(n5012), .B1(n4563), .B2(n1885), .ZN(n4539)
         );
  nd02d0 U3036 ( .A1(n2013), .A2(mprj_dat_o[7]), .ZN(n2635) );
  aoi22d1 U3037 ( .A1(n1886), .A2(n2635), .B1(n4567), .B2(n1885), .ZN(n4538)
         );
  nr02d0 U3038 ( .A1(count[0]), .A2(n1887), .ZN(n4537) );
  inv0d0 U3039 ( .I(request[1]), .ZN(n1897) );
  oai211d1 U3040 ( .C1(n1898), .C2(request[0]), .A(n1888), .B(n1897), .ZN(
        n1889) );
  oai211d1 U3041 ( .C1(request[0]), .C2(n1890), .A(n4881), .B(n1889), .ZN(
        n1896) );
  oai211d1 U3042 ( .C1(request[1]), .C2(request[0]), .A(n1891), .B(n1895), 
        .ZN(n1892) );
  nd12d0 U3043 ( .A1(n1896), .A2(n1892), .ZN(n1901) );
  oai21d1 U3044 ( .B1(n1896), .B2(n1895), .A(n1894), .ZN(n4517) );
  oai21d1 U3045 ( .B1(n1901), .B2(n1900), .A(n1899), .ZN(n4516) );
  nr02d0 U3046 ( .A1(n1937), .A2(n4575), .ZN(n1905) );
  oai21d1 U3047 ( .B1(gpioin5_i02), .B2(n1905), .A(n4881), .ZN(n1904) );
  aoi21d1 U3048 ( .B1(n1905), .B2(n4808), .A(n1904), .ZN(n4515) );
  oai21d1 U3049 ( .B1(gpioin5_pending_r), .B2(n1907), .A(n5301), .ZN(n1906) );
  aoi21d1 U3050 ( .B1(n1907), .B2(n4808), .A(n1906), .ZN(n4514) );
  inv0d0 U3051 ( .I(n4575), .ZN(n2647) );
  nd02d0 U3052 ( .A1(n2647), .A2(n1944), .ZN(n1909) );
  nd02d0 U3053 ( .A1(n4582), .A2(n5340), .ZN(n5000) );
  buffd1 U3054 ( .I(n5000), .Z(n4955) );
  nd03d0 U3055 ( .A1(n1909), .A2(gpioin4_i02), .A3(n5301), .ZN(n1908) );
  oai21d1 U3056 ( .B1(n1909), .B2(n4955), .A(n1908), .ZN(n4513) );
  oai21d1 U3057 ( .B1(n1911), .B2(n4955), .A(n1910), .ZN(n4512) );
  nd02d0 U3058 ( .A1(n2647), .A2(n1912), .ZN(n1914) );
  nd03d0 U3059 ( .A1(n1914), .A2(gpioin3_i02), .A3(n5956), .ZN(n1913) );
  oai21d1 U3060 ( .B1(n1914), .B2(n5000), .A(n1913), .ZN(n4511) );
  oai21d1 U3061 ( .B1(gpioin3_pending_r), .B2(n1916), .A(n5319), .ZN(n1915) );
  aoi21d1 U3062 ( .B1(n1916), .B2(n5290), .A(n1915), .ZN(n4510) );
  nr02d0 U3063 ( .A1(n4575), .A2(n1959), .ZN(n1918) );
  oai21d1 U3064 ( .B1(gpioin2_i02), .B2(n1918), .A(n5319), .ZN(n1917) );
  aoi21d1 U3065 ( .B1(n1918), .B2(n4808), .A(n1917), .ZN(n4509) );
  nr02d0 U3066 ( .A1(n1959), .A2(n2654), .ZN(n1920) );
  oai21d1 U3067 ( .B1(gpioin2_pending_r), .B2(n1920), .A(n5319), .ZN(n1919) );
  aoi21d1 U3068 ( .B1(n1920), .B2(n4808), .A(n1919), .ZN(n4508) );
  nr02d0 U3069 ( .A1(n4575), .A2(n1966), .ZN(n1922) );
  oai21d1 U3070 ( .B1(gpioin1_i02), .B2(n1922), .A(n5955), .ZN(n1921) );
  aoi21d1 U3071 ( .B1(n1922), .B2(n5290), .A(n1921), .ZN(n4507) );
  oai21d1 U3072 ( .B1(gpioin1_pending_r), .B2(n1924), .A(n5956), .ZN(n1923) );
  aoi21d1 U3073 ( .B1(n1924), .B2(n5290), .A(n1923), .ZN(n4506) );
  nr02d0 U3074 ( .A1(n4575), .A2(n1973), .ZN(n1926) );
  oai21d1 U3075 ( .B1(gpioin0_i02), .B2(n1926), .A(n4881), .ZN(n1925) );
  aoi21d1 U3076 ( .B1(n1926), .B2(n4808), .A(n1925), .ZN(n4505) );
  oai21d1 U3077 ( .B1(gpioin0_pending_r), .B2(n1928), .A(n5955), .ZN(n1927) );
  aoi21d1 U3078 ( .B1(n1928), .B2(n5290), .A(n1927), .ZN(n4504) );
  nd02d0 U3079 ( .A1(litespi_tx_mux_sel), .A2(\litespi_request[1] ), .ZN(n4846) );
  aoi211d1 U3080 ( .C1(mgmtsoc_litespimmap_burst_cs), .C2(n1930), .A(n1929), 
        .B(n4843), .ZN(n4847) );
  inv0d0 U3081 ( .I(n4847), .ZN(n1932) );
  oai21d1 U3082 ( .B1(litespi_tx_mux_sel), .B2(\litespi_request[1] ), .A(n5319), .ZN(n1931) );
  aoi21d1 U3083 ( .B1(n4846), .B2(n1932), .A(n1931), .ZN(n4503) );
  oaim21d1 U3084 ( .B1(gpioin5_pending_r), .B2(gpioin5_pending_re), .A(
        gpioin5_i01), .ZN(n1933) );
  oan211d1 U3085 ( .C1(n1934), .C2(gpioin5_gpioin5_trigger_d), .B(n1933), .A(
        n5100), .ZN(n4502) );
  nr02d0 U3086 ( .A1(n1937), .A2(n2334), .ZN(n1936) );
  oai21d1 U3087 ( .B1(csrbank18_edge0_w), .B2(n1936), .A(n5319), .ZN(n1935) );
  aoi21d1 U3088 ( .B1(n1936), .B2(n4808), .A(n1935), .ZN(n4501) );
  oai21d1 U3089 ( .B1(csrbank18_mode0_w), .B2(n1939), .A(n4881), .ZN(n1938) );
  aoi21d1 U3090 ( .B1(n1939), .B2(n4808), .A(n1938), .ZN(n4500) );
  oaim21d1 U3091 ( .B1(gpioin4_pending_r), .B2(gpioin4_pending_re), .A(
        gpioin4_i01), .ZN(n1940) );
  oan211d1 U3092 ( .C1(n1941), .C2(gpioin4_gpioin4_trigger_d), .B(n1940), .A(
        n4878), .ZN(n4499) );
  inv0d0 U3093 ( .I(n2334), .ZN(n2335) );
  nd02d0 U3094 ( .A1(n1944), .A2(n2335), .ZN(n1943) );
  oai21d1 U3095 ( .B1(n1943), .B2(n4955), .A(n1942), .ZN(n4498) );
  inv0d0 U3096 ( .I(n4959), .ZN(n5240) );
  nd02d0 U3097 ( .A1(n1944), .A2(n5240), .ZN(n1946) );
  oai21d1 U3098 ( .B1(n4582), .B2(n1946), .A(n5956), .ZN(n1945) );
  aoi21d1 U3099 ( .B1(n1947), .B2(n1946), .A(n1945), .ZN(n4497) );
  oaim21d1 U3100 ( .B1(gpioin3_pending_r), .B2(gpioin3_pending_re), .A(
        gpioin3_i01), .ZN(n1948) );
  oan211d1 U3101 ( .C1(n1949), .C2(gpioin3_gpioin3_trigger_d), .B(n1948), .A(
        sys_rst), .ZN(n4496) );
  nr02d0 U3102 ( .A1(n1952), .A2(n2334), .ZN(n1951) );
  oai21d1 U3103 ( .B1(csrbank16_edge0_w), .B2(n1951), .A(n5319), .ZN(n1950) );
  aoi21d1 U3104 ( .B1(n1951), .B2(n4808), .A(n1950), .ZN(n4495) );
  oai21d1 U3105 ( .B1(csrbank16_mode0_w), .B2(n1954), .A(n5340), .ZN(n1953) );
  aoi21d1 U3106 ( .B1(n1954), .B2(n4808), .A(n1953), .ZN(n4494) );
  inv0d0 U3107 ( .I(N6223), .ZN(n1956) );
  oaim21d1 U3108 ( .B1(gpioin2_pending_r), .B2(gpioin2_pending_re), .A(
        gpioin2_i01), .ZN(n1955) );
  oai22d1 U3109 ( .A1(gpioin2_gpioin2_trigger_d), .A2(n1956), .B1(sys_rst), 
        .B2(n1955), .ZN(n4493) );
  nr02d0 U3110 ( .A1(n1959), .A2(n2334), .ZN(n1958) );
  oai21d1 U3111 ( .B1(csrbank15_edge0_w), .B2(n1958), .A(n5319), .ZN(n1957) );
  aoi21d1 U3112 ( .B1(n1958), .B2(n4808), .A(n1957), .ZN(n4492) );
  nr02d0 U3113 ( .A1(n1959), .A2(n4959), .ZN(n1961) );
  oai21d1 U3114 ( .B1(csrbank15_mode0_w), .B2(n1961), .A(n5319), .ZN(n1960) );
  aoi21d1 U3115 ( .B1(n1961), .B2(n5290), .A(n1960), .ZN(n4491) );
  inv0d0 U3116 ( .I(N6215), .ZN(n1963) );
  oaim21d1 U3117 ( .B1(gpioin1_pending_r), .B2(gpioin1_pending_re), .A(
        gpioin1_i01), .ZN(n1962) );
  oai22d1 U3118 ( .A1(gpioin1_gpioin1_trigger_d), .A2(n1963), .B1(sys_rst), 
        .B2(n1962), .ZN(n4490) );
  nr02d0 U3119 ( .A1(n1966), .A2(n2334), .ZN(n1965) );
  oai21d1 U3120 ( .B1(csrbank14_edge0_w), .B2(n1965), .A(n5319), .ZN(n1964) );
  aoi21d1 U3121 ( .B1(n1965), .B2(n5290), .A(n1964), .ZN(n4489) );
  oai21d1 U3122 ( .B1(csrbank14_mode0_w), .B2(n1968), .A(n5319), .ZN(n1967) );
  aoi21d1 U3123 ( .B1(n1968), .B2(n5290), .A(n1967), .ZN(n4488) );
  inv0d0 U3124 ( .I(N6207), .ZN(n1970) );
  oaim21d1 U3125 ( .B1(gpioin0_pending_r), .B2(gpioin0_pending_re), .A(
        gpioin0_i01), .ZN(n1969) );
  oai22d1 U3126 ( .A1(gpioin0_gpioin0_trigger_d), .A2(n1970), .B1(n2516), .B2(
        n1969), .ZN(n4487) );
  oai21d1 U3127 ( .B1(csrbank13_edge0_w), .B2(n1972), .A(n5319), .ZN(n1971) );
  aoi21d1 U3128 ( .B1(n1972), .B2(n5290), .A(n1971), .ZN(n4486) );
  nr02d0 U3129 ( .A1(n1973), .A2(n4959), .ZN(n1975) );
  inv0d0 U3130 ( .I(n4582), .ZN(n2472) );
  oai21d1 U3131 ( .B1(csrbank13_mode0_w), .B2(n1975), .A(n5319), .ZN(n1974) );
  aoi21d1 U3132 ( .B1(n1975), .B2(n2472), .A(n1974), .ZN(n4485) );
  or02d0 U3133 ( .A1(n1976), .A2(n4811), .Z(n1981) );
  oai22d1 U3134 ( .A1(n4955), .A2(n1981), .B1(n1980), .B2(n1977), .ZN(n4484)
         );
  nd12d0 U3135 ( .A1(n4862), .A2(n5301), .ZN(n2653) );
  oai22d1 U3136 ( .A1(n2653), .A2(n1981), .B1(n1980), .B2(n1978), .ZN(n4483)
         );
  oai22d1 U3137 ( .A1(n2298), .A2(n1981), .B1(n1980), .B2(n1979), .ZN(n4482)
         );
  nd03d0 U3138 ( .A1(n1984), .A2(spi_enabled), .A3(n5301), .ZN(n1983) );
  oai21d1 U3139 ( .B1(n1984), .B2(n4955), .A(n1983), .ZN(n4481) );
  inv0d0 U3140 ( .I(n134), .ZN(n1986) );
  nd02d1 U3141 ( .A1(n5955), .A2(n1989), .ZN(n2015) );
  aoi22d1 U3142 ( .A1(n1986), .A2(n1989), .B1(n4955), .B2(n2015), .ZN(n4480)
         );
  inv0d0 U3143 ( .I(n133), .ZN(n1987) );
  aoi22d1 U3144 ( .A1(n1987), .A2(n1989), .B1(n2015), .B2(n2653), .ZN(n4479)
         );
  inv0d0 U3145 ( .I(n132), .ZN(n1988) );
  aoi22d1 U3146 ( .A1(n1988), .A2(n1989), .B1(n2015), .B2(n2298), .ZN(n4478)
         );
  inv0d0 U3147 ( .I(n131), .ZN(n1990) );
  or02d1 U3148 ( .A1(n1989), .A2(n5111), .Z(n2020) );
  oai22d1 U3149 ( .A1(n1990), .A2(n2015), .B1(n2625), .B2(n2020), .ZN(n4477)
         );
  inv0d0 U3150 ( .I(n130), .ZN(n1991) );
  buffd1 U3151 ( .I(n2020), .Z(n2023) );
  oai22d1 U3152 ( .A1(n1991), .A2(n2015), .B1(n4866), .B2(n2023), .ZN(n4476)
         );
  inv0d0 U3153 ( .I(n129), .ZN(n1992) );
  buffd1 U3154 ( .I(n2015), .Z(n2024) );
  buffd1 U3155 ( .I(n2640), .Z(n5248) );
  oai22d1 U3156 ( .A1(n1992), .A2(n2024), .B1(n5248), .B2(n2023), .ZN(n4475)
         );
  inv0d0 U3157 ( .I(n128), .ZN(n1993) );
  buffd1 U3158 ( .I(n2641), .Z(n5249) );
  oai22d1 U3159 ( .A1(n1993), .A2(n2015), .B1(n5249), .B2(n2023), .ZN(n4474)
         );
  inv0d0 U3160 ( .I(n127), .ZN(n1994) );
  buffd1 U3161 ( .I(n2635), .Z(n3071) );
  oai22d1 U3162 ( .A1(n1994), .A2(n2015), .B1(n3071), .B2(n2023), .ZN(n4473)
         );
  inv0d0 U3163 ( .I(n126), .ZN(n1995) );
  nd02d1 U3164 ( .A1(n2022), .A2(mprj_dat_o[8]), .ZN(n4783) );
  inv0d0 U3165 ( .I(n4783), .ZN(n2035) );
  inv0d0 U3166 ( .I(n2035), .ZN(n5015) );
  oai22d1 U3167 ( .A1(n1995), .A2(n2015), .B1(n2023), .B2(n5015), .ZN(n4472)
         );
  inv0d0 U3168 ( .I(n125), .ZN(n1996) );
  nd02d1 U3169 ( .A1(n2022), .A2(mprj_dat_o[9]), .ZN(n4593) );
  inv0d0 U3170 ( .I(n4593), .ZN(n2077) );
  inv0d0 U3171 ( .I(n2077), .ZN(n5017) );
  oai22d1 U3172 ( .A1(n1996), .A2(n2024), .B1(n2023), .B2(n5017), .ZN(n4471)
         );
  inv0d0 U3173 ( .I(n124), .ZN(n1997) );
  nd02d1 U3174 ( .A1(n2022), .A2(mprj_dat_o[10]), .ZN(n4595) );
  inv0d0 U3175 ( .I(n4595), .ZN(n2079) );
  inv0d0 U3176 ( .I(n2079), .ZN(n5019) );
  oai22d1 U3177 ( .A1(n1997), .A2(n2015), .B1(n2023), .B2(n5019), .ZN(n4470)
         );
  inv0d0 U3178 ( .I(n123), .ZN(n1998) );
  nd02d1 U3179 ( .A1(n2022), .A2(mprj_dat_o[11]), .ZN(n4787) );
  inv0d0 U3180 ( .I(n4787), .ZN(n2039) );
  oai22d1 U3181 ( .A1(n1998), .A2(n2024), .B1(n2023), .B2(n4787), .ZN(n4469)
         );
  inv0d0 U3182 ( .I(n122), .ZN(n1999) );
  nd02d1 U3183 ( .A1(n2022), .A2(mprj_dat_o[12]), .ZN(n4598) );
  inv0d0 U3184 ( .I(n4598), .ZN(n2082) );
  inv0d0 U3185 ( .I(n2082), .ZN(n5022) );
  oai22d1 U3186 ( .A1(n1999), .A2(n2024), .B1(n2023), .B2(n5022), .ZN(n4468)
         );
  inv0d0 U3187 ( .I(n121), .ZN(n2000) );
  nd02d1 U3188 ( .A1(n2022), .A2(mprj_dat_o[13]), .ZN(n4790) );
  inv0d0 U3189 ( .I(n4790), .ZN(n2042) );
  inv0d0 U3190 ( .I(n2042), .ZN(n5024) );
  oai22d1 U3191 ( .A1(n2000), .A2(n2024), .B1(n2023), .B2(n5024), .ZN(n4467)
         );
  inv0d0 U3192 ( .I(n120), .ZN(n2001) );
  nd02d1 U3193 ( .A1(n2022), .A2(mprj_dat_o[14]), .ZN(n4601) );
  inv0d0 U3194 ( .I(n4601), .ZN(n2085) );
  inv0d0 U3195 ( .I(n2085), .ZN(n5026) );
  oai22d1 U3196 ( .A1(n2001), .A2(n2015), .B1(n2020), .B2(n5026), .ZN(n4466)
         );
  inv0d0 U3197 ( .I(n119), .ZN(n2002) );
  nd02d1 U3198 ( .A1(n2022), .A2(mprj_dat_o[15]), .ZN(n4793) );
  inv0d0 U3199 ( .I(n4793), .ZN(n2045) );
  inv0d0 U3200 ( .I(n2045), .ZN(n5028) );
  oai22d1 U3201 ( .A1(n2002), .A2(n2015), .B1(n2020), .B2(n5028), .ZN(n4465)
         );
  inv0d0 U3202 ( .I(n118), .ZN(n2004) );
  nd02d1 U3203 ( .A1(n2022), .A2(mprj_dat_o[16]), .ZN(n2003) );
  oai22d1 U3204 ( .A1(n2004), .A2(n2024), .B1(n2023), .B2(n2003), .ZN(n4464)
         );
  inv0d0 U3205 ( .I(n117), .ZN(n2005) );
  nd02d1 U3206 ( .A1(n2022), .A2(mprj_dat_o[17]), .ZN(n5259) );
  oai22d1 U3207 ( .A1(n2005), .A2(n2024), .B1(n2023), .B2(n5259), .ZN(n4463)
         );
  inv0d0 U3208 ( .I(n116), .ZN(n2006) );
  nd02d1 U3209 ( .A1(n2013), .A2(mprj_dat_o[18]), .ZN(n5260) );
  oai22d1 U3210 ( .A1(n2006), .A2(n2015), .B1(n2023), .B2(n5260), .ZN(n4462)
         );
  inv0d0 U3211 ( .I(n115), .ZN(n2007) );
  nd02d1 U3212 ( .A1(n2022), .A2(mprj_dat_o[19]), .ZN(n5262) );
  oai22d1 U3213 ( .A1(n2007), .A2(n2015), .B1(n2023), .B2(n5262), .ZN(n4461)
         );
  inv0d0 U3214 ( .I(n114), .ZN(n2008) );
  nd02d1 U3215 ( .A1(n2013), .A2(mprj_dat_o[20]), .ZN(n5263) );
  oai22d1 U3216 ( .A1(n2008), .A2(n2024), .B1(n2020), .B2(n5263), .ZN(n4460)
         );
  inv0d0 U3217 ( .I(n113), .ZN(n2009) );
  nd02d1 U3218 ( .A1(n2022), .A2(mprj_dat_o[21]), .ZN(n5264) );
  oai22d1 U3219 ( .A1(n2009), .A2(n2024), .B1(n2020), .B2(n5264), .ZN(n4459)
         );
  inv0d0 U3220 ( .I(n112), .ZN(n2010) );
  nd02d1 U3221 ( .A1(n2022), .A2(mprj_dat_o[22]), .ZN(n5266) );
  oai22d1 U3222 ( .A1(n2010), .A2(n2024), .B1(n2023), .B2(n5266), .ZN(n4458)
         );
  inv0d0 U3223 ( .I(n111), .ZN(n2011) );
  nd02d1 U3224 ( .A1(n2013), .A2(mprj_dat_o[23]), .ZN(n5268) );
  oai22d1 U3225 ( .A1(n2011), .A2(n2024), .B1(n2023), .B2(n5268), .ZN(n4457)
         );
  inv0d0 U3226 ( .I(n110), .ZN(n2012) );
  nd02d1 U3227 ( .A1(n2013), .A2(mprj_dat_o[24]), .ZN(n5270) );
  oai22d1 U3228 ( .A1(n2012), .A2(n2024), .B1(n2020), .B2(n5270), .ZN(n4456)
         );
  inv0d0 U3229 ( .I(n109), .ZN(n2014) );
  nd02d1 U3230 ( .A1(n2013), .A2(mprj_dat_o[25]), .ZN(n5271) );
  oai22d1 U3231 ( .A1(n2014), .A2(n2015), .B1(n2020), .B2(n5271), .ZN(n4455)
         );
  inv0d0 U3232 ( .I(n108), .ZN(n2016) );
  nd02d1 U3233 ( .A1(n2022), .A2(mprj_dat_o[26]), .ZN(n5273) );
  oai22d1 U3234 ( .A1(n2016), .A2(n2015), .B1(n2020), .B2(n5273), .ZN(n4454)
         );
  inv0d0 U3235 ( .I(n107), .ZN(n2017) );
  nd02d1 U3236 ( .A1(n2022), .A2(mprj_dat_o[27]), .ZN(n5275) );
  oai22d1 U3237 ( .A1(n2017), .A2(n2024), .B1(n2020), .B2(n5275), .ZN(n4453)
         );
  inv0d0 U3238 ( .I(n106), .ZN(n2018) );
  nd02d1 U3239 ( .A1(n2022), .A2(mprj_dat_o[28]), .ZN(n5276) );
  oai22d1 U3240 ( .A1(n2018), .A2(n2024), .B1(n2020), .B2(n5276), .ZN(n4452)
         );
  inv0d0 U3241 ( .I(n105), .ZN(n2019) );
  nd02d1 U3242 ( .A1(n2022), .A2(mprj_dat_o[29]), .ZN(n5280) );
  oai22d1 U3243 ( .A1(n2019), .A2(n2024), .B1(n2020), .B2(n5280), .ZN(n4451)
         );
  inv0d0 U3244 ( .I(n104), .ZN(n2021) );
  nd02d1 U3245 ( .A1(n2022), .A2(mprj_dat_o[30]), .ZN(n5283) );
  oai22d1 U3246 ( .A1(n2021), .A2(n2024), .B1(n2020), .B2(n5283), .ZN(n4450)
         );
  inv0d0 U3247 ( .I(n103), .ZN(n2025) );
  nd02d1 U3248 ( .A1(n2022), .A2(mprj_dat_o[31]), .ZN(n5287) );
  oai22d1 U3249 ( .A1(n2025), .A2(n2024), .B1(n2023), .B2(n5287), .ZN(n4449)
         );
  inv0d0 U3250 ( .I(n102), .ZN(n2027) );
  oaim21d1 U3251 ( .B1(n4683), .B2(n2026), .A(n5340), .ZN(n2057) );
  inv0d0 U3252 ( .I(n4957), .ZN(n4580) );
  nd02d1 U3253 ( .A1(n2026), .A2(n4580), .ZN(n2064) );
  buffd1 U3254 ( .I(n2064), .Z(n2053) );
  oai22d1 U3255 ( .A1(n2027), .A2(n2057), .B1(n5290), .B2(n2053), .ZN(n4448)
         );
  inv0d0 U3256 ( .I(n101), .ZN(n2028) );
  oai22d1 U3257 ( .A1(n2028), .A2(n2057), .B1(n4862), .B2(n2053), .ZN(n4447)
         );
  inv0d0 U3258 ( .I(n100), .ZN(n2029) );
  oai22d1 U3259 ( .A1(n2029), .A2(n2057), .B1(n5004), .B2(n2053), .ZN(n4446)
         );
  inv0d0 U3260 ( .I(n99), .ZN(n2030) );
  buffd1 U3261 ( .I(n2625), .Z(n5246) );
  oai22d1 U3262 ( .A1(n2030), .A2(n2057), .B1(n5246), .B2(n2053), .ZN(n4445)
         );
  inv0d0 U3263 ( .I(n98), .ZN(n2031) );
  buffd1 U3264 ( .I(n2057), .Z(n2065) );
  buffd1 U3265 ( .I(n4866), .Z(n5247) );
  oai22d1 U3266 ( .A1(n2031), .A2(n2065), .B1(n5247), .B2(n2053), .ZN(n4444)
         );
  inv0d0 U3267 ( .I(n97), .ZN(n2032) );
  oai22d1 U3268 ( .A1(n2032), .A2(n2057), .B1(n5248), .B2(n2053), .ZN(n4443)
         );
  inv0d0 U3269 ( .I(n96), .ZN(n2033) );
  oai22d1 U3270 ( .A1(n2033), .A2(n2057), .B1(n5249), .B2(n2053), .ZN(n4442)
         );
  inv0d0 U3271 ( .I(n95), .ZN(n2034) );
  oai22d1 U3272 ( .A1(n2034), .A2(n2057), .B1(n3071), .B2(n2053), .ZN(n4441)
         );
  inv0d0 U3273 ( .I(n94), .ZN(n2036) );
  oai22d1 U3274 ( .A1(n2036), .A2(n2065), .B1(n4783), .B2(n2053), .ZN(n4440)
         );
  inv0d0 U3275 ( .I(n93), .ZN(n2037) );
  oai22d1 U3276 ( .A1(n2037), .A2(n2065), .B1(n5017), .B2(n2053), .ZN(n4439)
         );
  inv0d0 U3277 ( .I(n92), .ZN(n2038) );
  oai22d1 U3278 ( .A1(n2038), .A2(n2065), .B1(n5019), .B2(n2064), .ZN(n4438)
         );
  inv0d0 U3279 ( .I(n91), .ZN(n2040) );
  inv0d0 U3280 ( .I(n2039), .ZN(n5254) );
  oai22d1 U3281 ( .A1(n2040), .A2(n2065), .B1(n5254), .B2(n2064), .ZN(n4437)
         );
  inv0d0 U3282 ( .I(n90), .ZN(n2041) );
  oai22d1 U3283 ( .A1(n2041), .A2(n2065), .B1(n5022), .B2(n2053), .ZN(n4436)
         );
  inv0d0 U3284 ( .I(n89), .ZN(n2043) );
  oai22d1 U3285 ( .A1(n2043), .A2(n2065), .B1(n4790), .B2(n2064), .ZN(n4435)
         );
  inv0d0 U3286 ( .I(n88), .ZN(n2044) );
  oai22d1 U3287 ( .A1(n2044), .A2(n2065), .B1(n5026), .B2(n2053), .ZN(n4434)
         );
  inv0d0 U3288 ( .I(n87), .ZN(n2046) );
  oai22d1 U3289 ( .A1(n2046), .A2(n2057), .B1(n4793), .B2(n2053), .ZN(n4433)
         );
  inv0d0 U3290 ( .I(n86), .ZN(n2047) );
  oai22d1 U3291 ( .A1(n2047), .A2(n2057), .B1(n2003), .B2(n2053), .ZN(n4432)
         );
  inv0d0 U3292 ( .I(n85), .ZN(n2048) );
  oai22d1 U3293 ( .A1(n2048), .A2(n2057), .B1(n5259), .B2(n2064), .ZN(n4431)
         );
  inv0d0 U3294 ( .I(n84), .ZN(n2049) );
  oai22d1 U3295 ( .A1(n2049), .A2(n2065), .B1(n5260), .B2(n2064), .ZN(n4430)
         );
  inv0d0 U3296 ( .I(n83), .ZN(n2050) );
  oai22d1 U3297 ( .A1(n2050), .A2(n2057), .B1(n5262), .B2(n2053), .ZN(n4429)
         );
  inv0d0 U3298 ( .I(n82), .ZN(n2051) );
  oai22d1 U3299 ( .A1(n2051), .A2(n2057), .B1(n5263), .B2(n2064), .ZN(n4428)
         );
  inv0d0 U3300 ( .I(n81), .ZN(n2052) );
  oai22d1 U3301 ( .A1(n2052), .A2(n2057), .B1(n5264), .B2(n2053), .ZN(n4427)
         );
  inv0d0 U3302 ( .I(n80), .ZN(n2054) );
  oai22d1 U3303 ( .A1(n2054), .A2(n2057), .B1(n5266), .B2(n2053), .ZN(n4426)
         );
  inv0d0 U3304 ( .I(n79), .ZN(n2055) );
  oai22d1 U3305 ( .A1(n2055), .A2(n2057), .B1(n5268), .B2(n2064), .ZN(n4425)
         );
  inv0d0 U3306 ( .I(n78), .ZN(n2056) );
  oai22d1 U3307 ( .A1(n2056), .A2(n2065), .B1(n5270), .B2(n2064), .ZN(n4424)
         );
  inv0d0 U3308 ( .I(n77), .ZN(n2058) );
  oai22d1 U3309 ( .A1(n2058), .A2(n2057), .B1(n5271), .B2(n2064), .ZN(n4423)
         );
  inv0d0 U3310 ( .I(n76), .ZN(n2059) );
  oai22d1 U3311 ( .A1(n2059), .A2(n2065), .B1(n5273), .B2(n2064), .ZN(n4422)
         );
  inv0d0 U3312 ( .I(n75), .ZN(n2060) );
  oai22d1 U3313 ( .A1(n2060), .A2(n2065), .B1(n5275), .B2(n2064), .ZN(n4421)
         );
  inv0d0 U3314 ( .I(n74), .ZN(n2061) );
  oai22d1 U3315 ( .A1(n2061), .A2(n2065), .B1(n5276), .B2(n2064), .ZN(n4420)
         );
  inv0d0 U3316 ( .I(n73), .ZN(n2062) );
  oai22d1 U3317 ( .A1(n2062), .A2(n2065), .B1(n5280), .B2(n2064), .ZN(n4419)
         );
  inv0d0 U3318 ( .I(n72), .ZN(n2063) );
  oai22d1 U3319 ( .A1(n2063), .A2(n2065), .B1(n5283), .B2(n2064), .ZN(n4418)
         );
  inv0d0 U3320 ( .I(n71), .ZN(n2066) );
  oai22d1 U3321 ( .A1(n2066), .A2(n2065), .B1(n5287), .B2(n2064), .ZN(n4417)
         );
  inv0d0 U3322 ( .I(n70), .ZN(n2068) );
  nd02d1 U3323 ( .A1(n2067), .A2(n4580), .ZN(n2105) );
  buffd1 U3324 ( .I(n2105), .Z(n2103) );
  nd02d1 U3325 ( .A1(n5288), .A2(n2103), .ZN(n2098) );
  oai22d1 U3326 ( .A1(n2068), .A2(n2098), .B1(n4808), .B2(n2103), .ZN(n4416)
         );
  inv0d0 U3327 ( .I(n69), .ZN(n2069) );
  oai22d1 U3328 ( .A1(n2069), .A2(n2098), .B1(n2639), .B2(n2103), .ZN(n4415)
         );
  inv0d0 U3329 ( .I(n68), .ZN(n2070) );
  oai22d1 U3330 ( .A1(n2070), .A2(n2098), .B1(n5004), .B2(n2103), .ZN(n4414)
         );
  inv0d0 U3331 ( .I(n67), .ZN(n2071) );
  oai22d1 U3332 ( .A1(n2071), .A2(n2098), .B1(n5246), .B2(n2103), .ZN(n4413)
         );
  inv0d0 U3333 ( .I(n66), .ZN(n2072) );
  buffd1 U3334 ( .I(n2098), .Z(n2106) );
  oai22d1 U3335 ( .A1(n2072), .A2(n2106), .B1(n5247), .B2(n2103), .ZN(n4412)
         );
  inv0d0 U3336 ( .I(n65), .ZN(n2073) );
  oai22d1 U3337 ( .A1(n2073), .A2(n2098), .B1(n5248), .B2(n2103), .ZN(n4411)
         );
  inv0d0 U3338 ( .I(n64), .ZN(n2074) );
  oai22d1 U3339 ( .A1(n2074), .A2(n2098), .B1(n5249), .B2(n2103), .ZN(n4410)
         );
  inv0d0 U3340 ( .I(n63), .ZN(n2075) );
  oai22d1 U3341 ( .A1(n2075), .A2(n2098), .B1(n3071), .B2(n2105), .ZN(n4409)
         );
  inv0d0 U3342 ( .I(n62), .ZN(n2076) );
  oai22d1 U3343 ( .A1(n2076), .A2(n2098), .B1(n4783), .B2(n2105), .ZN(n4408)
         );
  inv0d0 U3344 ( .I(n61), .ZN(n2078) );
  oai22d1 U3345 ( .A1(n2078), .A2(n2106), .B1(n4593), .B2(n2103), .ZN(n4407)
         );
  inv0d0 U3346 ( .I(n60), .ZN(n2080) );
  oai22d1 U3347 ( .A1(n2080), .A2(n2098), .B1(n4595), .B2(n2105), .ZN(n4406)
         );
  inv0d0 U3348 ( .I(n59), .ZN(n2081) );
  oai22d1 U3349 ( .A1(n2081), .A2(n2098), .B1(n5254), .B2(n2105), .ZN(n4405)
         );
  inv0d0 U3350 ( .I(n58), .ZN(n2083) );
  oai22d1 U3351 ( .A1(n2083), .A2(n2106), .B1(n4598), .B2(n2103), .ZN(n4404)
         );
  inv0d0 U3352 ( .I(n57), .ZN(n2084) );
  oai22d1 U3353 ( .A1(n2084), .A2(n2106), .B1(n4790), .B2(n2103), .ZN(n4403)
         );
  inv0d0 U3354 ( .I(n56), .ZN(n2086) );
  oai22d1 U3355 ( .A1(n2086), .A2(n2098), .B1(n4601), .B2(n2105), .ZN(n4402)
         );
  inv0d0 U3356 ( .I(n55), .ZN(n2087) );
  oai22d1 U3357 ( .A1(n2087), .A2(n2098), .B1(n4793), .B2(n2105), .ZN(n4401)
         );
  inv0d0 U3358 ( .I(n54), .ZN(n2088) );
  oai22d1 U3359 ( .A1(n2088), .A2(n2106), .B1(n2003), .B2(n2105), .ZN(n4400)
         );
  inv0d0 U3360 ( .I(n53), .ZN(n2089) );
  oai22d1 U3361 ( .A1(n2089), .A2(n2106), .B1(n5259), .B2(n2105), .ZN(n4399)
         );
  inv0d0 U3362 ( .I(n52), .ZN(n2090) );
  oai22d1 U3363 ( .A1(n2090), .A2(n2106), .B1(n5260), .B2(n2105), .ZN(n4398)
         );
  inv0d0 U3364 ( .I(n51), .ZN(n2091) );
  oai22d1 U3365 ( .A1(n2091), .A2(n2106), .B1(n5262), .B2(n2105), .ZN(n4397)
         );
  inv0d0 U3366 ( .I(n50), .ZN(n2092) );
  oai22d1 U3367 ( .A1(n2092), .A2(n2106), .B1(n5263), .B2(n2105), .ZN(n4396)
         );
  inv0d0 U3368 ( .I(n49), .ZN(n2093) );
  oai22d1 U3369 ( .A1(n2093), .A2(n2106), .B1(n5264), .B2(n2103), .ZN(n4395)
         );
  inv0d0 U3370 ( .I(n48), .ZN(n2094) );
  oai22d1 U3371 ( .A1(n2094), .A2(n2098), .B1(n5266), .B2(n2103), .ZN(n4394)
         );
  inv0d0 U3372 ( .I(n47), .ZN(n2095) );
  oai22d1 U3373 ( .A1(n2095), .A2(n2106), .B1(n5268), .B2(n2103), .ZN(n4393)
         );
  inv0d0 U3374 ( .I(n46), .ZN(n2096) );
  oai22d1 U3375 ( .A1(n2096), .A2(n2098), .B1(n5270), .B2(n2105), .ZN(n4392)
         );
  inv0d0 U3376 ( .I(n45), .ZN(n2097) );
  oai22d1 U3377 ( .A1(n2097), .A2(n2106), .B1(n5271), .B2(n2103), .ZN(n4391)
         );
  inv0d0 U3378 ( .I(n44), .ZN(n2099) );
  oai22d1 U3379 ( .A1(n2099), .A2(n2098), .B1(n5273), .B2(n2105), .ZN(n4390)
         );
  inv0d0 U3380 ( .I(n43), .ZN(n2100) );
  oai22d1 U3381 ( .A1(n2100), .A2(n2106), .B1(n5275), .B2(n2103), .ZN(n4389)
         );
  inv0d0 U3382 ( .I(n42), .ZN(n2101) );
  oai22d1 U3383 ( .A1(n2101), .A2(n2106), .B1(n5276), .B2(n2105), .ZN(n4388)
         );
  inv0d0 U3384 ( .I(n41), .ZN(n2102) );
  oai22d1 U3385 ( .A1(n2102), .A2(n2106), .B1(n5280), .B2(n2105), .ZN(n4387)
         );
  inv0d0 U3386 ( .I(n40), .ZN(n2104) );
  oai22d1 U3387 ( .A1(n2104), .A2(n2106), .B1(n5283), .B2(n2103), .ZN(n4386)
         );
  inv0d0 U3388 ( .I(n39), .ZN(n2107) );
  oai22d1 U3389 ( .A1(n2107), .A2(n2106), .B1(n5287), .B2(n2105), .ZN(n4385)
         );
  inv0d0 U3390 ( .I(n38), .ZN(n2109) );
  nd02d1 U3391 ( .A1(n2108), .A2(n4580), .ZN(n2131) );
  nd02d1 U3392 ( .A1(n5288), .A2(n2131), .ZN(n2135) );
  buffd1 U3393 ( .I(n2131), .Z(n2142) );
  oai22d1 U3394 ( .A1(n2109), .A2(n2135), .B1(n4808), .B2(n2142), .ZN(n4384)
         );
  inv0d0 U3395 ( .I(n37), .ZN(n2110) );
  oai22d1 U3396 ( .A1(n2110), .A2(n2135), .B1(n5294), .B2(n2142), .ZN(n4383)
         );
  inv0d0 U3397 ( .I(n36), .ZN(n2111) );
  oai22d1 U3398 ( .A1(n2111), .A2(n2135), .B1(n5004), .B2(n2142), .ZN(n4382)
         );
  inv0d0 U3399 ( .I(n35), .ZN(n2112) );
  oai22d1 U3400 ( .A1(n2112), .A2(n2135), .B1(n5246), .B2(n2142), .ZN(n4381)
         );
  inv0d0 U3401 ( .I(n34), .ZN(n2113) );
  buffd1 U3402 ( .I(n2135), .Z(n2143) );
  oai22d1 U3403 ( .A1(n2113), .A2(n2143), .B1(n5247), .B2(n2142), .ZN(n4380)
         );
  inv0d0 U3404 ( .I(n33), .ZN(n2114) );
  oai22d1 U3405 ( .A1(n2114), .A2(n2135), .B1(n5248), .B2(n2131), .ZN(n4379)
         );
  inv0d0 U3406 ( .I(n32), .ZN(n2115) );
  oai22d1 U3407 ( .A1(n2115), .A2(n2143), .B1(n5249), .B2(n2131), .ZN(n4378)
         );
  inv0d0 U3408 ( .I(n31), .ZN(n2116) );
  buffd1 U3409 ( .I(n2635), .Z(n5251) );
  oai22d1 U3410 ( .A1(n2116), .A2(n2135), .B1(n5251), .B2(n2142), .ZN(n4377)
         );
  inv0d0 U3411 ( .I(n30), .ZN(n2117) );
  oai22d1 U3412 ( .A1(n2117), .A2(n2135), .B1(n5015), .B2(n2131), .ZN(n4376)
         );
  inv0d0 U3413 ( .I(n29), .ZN(n2118) );
  oai22d1 U3414 ( .A1(n2118), .A2(n2143), .B1(n5017), .B2(n2131), .ZN(n4375)
         );
  inv0d0 U3415 ( .I(n28), .ZN(n2119) );
  oai22d1 U3416 ( .A1(n2119), .A2(n2143), .B1(n5019), .B2(n2131), .ZN(n4374)
         );
  inv0d0 U3417 ( .I(n27), .ZN(n2120) );
  oai22d1 U3418 ( .A1(n2120), .A2(n2143), .B1(n4787), .B2(n2131), .ZN(n4373)
         );
  inv0d0 U3419 ( .I(n26), .ZN(n2121) );
  oai22d1 U3420 ( .A1(n2121), .A2(n2143), .B1(n5022), .B2(n2142), .ZN(n4372)
         );
  inv0d0 U3421 ( .I(n25), .ZN(n2122) );
  oai22d1 U3422 ( .A1(n2122), .A2(n2143), .B1(n5024), .B2(n2131), .ZN(n4371)
         );
  inv0d0 U3423 ( .I(n24), .ZN(n2123) );
  oai22d1 U3424 ( .A1(n2123), .A2(n2143), .B1(n5026), .B2(n2131), .ZN(n4370)
         );
  inv0d0 U3425 ( .I(n23), .ZN(n2124) );
  oai22d1 U3426 ( .A1(n2124), .A2(n2143), .B1(n5028), .B2(n2131), .ZN(n4369)
         );
  inv0d0 U3427 ( .I(n22), .ZN(n2125) );
  oai22d1 U3428 ( .A1(n2125), .A2(n2135), .B1(n2003), .B2(n2131), .ZN(n4368)
         );
  inv0d0 U3429 ( .I(n21), .ZN(n2126) );
  oai22d1 U3430 ( .A1(n2126), .A2(n2135), .B1(n5259), .B2(n2131), .ZN(n4367)
         );
  inv0d0 U3431 ( .I(n20), .ZN(n2127) );
  oai22d1 U3432 ( .A1(n2127), .A2(n2135), .B1(n5260), .B2(n2142), .ZN(n4366)
         );
  inv0d0 U3433 ( .I(n19), .ZN(n2128) );
  oai22d1 U3434 ( .A1(n2128), .A2(n2135), .B1(n5262), .B2(n2131), .ZN(n4365)
         );
  inv0d0 U3435 ( .I(n18), .ZN(n2129) );
  oai22d1 U3436 ( .A1(n2129), .A2(n2135), .B1(n5263), .B2(n2131), .ZN(n4364)
         );
  inv0d0 U3437 ( .I(n17), .ZN(n2130) );
  oai22d1 U3438 ( .A1(n2130), .A2(n2143), .B1(n5264), .B2(n2131), .ZN(n4363)
         );
  inv0d0 U3439 ( .I(n16), .ZN(n2132) );
  oai22d1 U3440 ( .A1(n2132), .A2(n2135), .B1(n5266), .B2(n2131), .ZN(n4362)
         );
  inv0d0 U3441 ( .I(n15), .ZN(n2133) );
  oai22d1 U3442 ( .A1(n2133), .A2(n2143), .B1(n5268), .B2(n2142), .ZN(n4361)
         );
  inv0d0 U3443 ( .I(n14), .ZN(n2134) );
  oai22d1 U3444 ( .A1(n2134), .A2(n2135), .B1(n5270), .B2(n2142), .ZN(n4360)
         );
  inv0d0 U3445 ( .I(n13), .ZN(n2136) );
  oai22d1 U3446 ( .A1(n2136), .A2(n2135), .B1(n5271), .B2(n2142), .ZN(n4359)
         );
  inv0d0 U3447 ( .I(n12), .ZN(n2137) );
  oai22d1 U3448 ( .A1(n2137), .A2(n2143), .B1(n5273), .B2(n2142), .ZN(n4358)
         );
  inv0d0 U3449 ( .I(n11), .ZN(n2138) );
  oai22d1 U3450 ( .A1(n2138), .A2(n2143), .B1(n5275), .B2(n2142), .ZN(n4357)
         );
  inv0d0 U3451 ( .I(n10), .ZN(n2139) );
  oai22d1 U3452 ( .A1(n2139), .A2(n2143), .B1(n5276), .B2(n2142), .ZN(n4356)
         );
  inv0d0 U3453 ( .I(n9), .ZN(n2140) );
  oai22d1 U3454 ( .A1(n2140), .A2(n2143), .B1(n5280), .B2(n2142), .ZN(n4355)
         );
  inv0d0 U3455 ( .I(n8), .ZN(n2141) );
  oai22d1 U3456 ( .A1(n2141), .A2(n2143), .B1(n5283), .B2(n2142), .ZN(n4354)
         );
  inv0d0 U3457 ( .I(n7), .ZN(n2144) );
  oai22d1 U3458 ( .A1(n2144), .A2(n2143), .B1(n5287), .B2(n2142), .ZN(n4353)
         );
  inv0d0 U3459 ( .I(csrbank6_oe0_w[0]), .ZN(n2145) );
  oaim21d1 U3460 ( .B1(n4683), .B2(n2148), .A(n4881), .ZN(n2181) );
  buffd1 U3461 ( .I(n2181), .Z(n2178) );
  nd02d0 U3462 ( .A1(n4683), .A2(n2148), .ZN(n2146) );
  oai22d1 U3463 ( .A1(n2145), .A2(n2178), .B1(n4955), .B2(n2146), .ZN(n4352)
         );
  inv0d0 U3464 ( .I(csrbank6_oe0_w[1]), .ZN(n2147) );
  aoi22d1 U3465 ( .A1(n2147), .A2(n2146), .B1(n2653), .B2(n2181), .ZN(n4351)
         );
  inv0d0 U3466 ( .I(csrbank6_oe0_w[2]), .ZN(n2149) );
  buffd3 U3467 ( .I(n2166), .Z(n2180) );
  oai22d1 U3468 ( .A1(n2149), .A2(n2178), .B1(n5004), .B2(n2180), .ZN(n4350)
         );
  inv0d0 U3469 ( .I(csrbank6_oe0_w[3]), .ZN(n2150) );
  oai22d1 U3470 ( .A1(n2150), .A2(n2178), .B1(n5246), .B2(n2180), .ZN(n4349)
         );
  inv0d0 U3471 ( .I(csrbank6_oe0_w[4]), .ZN(n2151) );
  oai22d1 U3472 ( .A1(n2151), .A2(n2178), .B1(n5247), .B2(n2180), .ZN(n4348)
         );
  inv0d0 U3473 ( .I(csrbank6_oe0_w[5]), .ZN(n2152) );
  oai22d1 U3474 ( .A1(n2152), .A2(n2178), .B1(n5248), .B2(n2180), .ZN(n4347)
         );
  inv0d0 U3475 ( .I(csrbank6_oe0_w[6]), .ZN(n2153) );
  oai22d1 U3476 ( .A1(n2153), .A2(n2178), .B1(n5249), .B2(n2180), .ZN(n4346)
         );
  inv0d0 U3477 ( .I(csrbank6_oe0_w[7]), .ZN(n2154) );
  oai22d1 U3478 ( .A1(n2154), .A2(n2181), .B1(n2635), .B2(n2180), .ZN(n4345)
         );
  inv0d0 U3479 ( .I(csrbank6_oe0_w[8]), .ZN(n2155) );
  oai22d1 U3480 ( .A1(n2155), .A2(n2181), .B1(n5015), .B2(n2180), .ZN(n4344)
         );
  inv0d0 U3481 ( .I(csrbank6_oe0_w[9]), .ZN(n2156) );
  oai22d1 U3482 ( .A1(n2156), .A2(n2178), .B1(n4593), .B2(n2180), .ZN(n4343)
         );
  inv0d0 U3483 ( .I(csrbank6_oe0_w[10]), .ZN(n2157) );
  oai22d1 U3484 ( .A1(n2157), .A2(n2178), .B1(n4595), .B2(n2180), .ZN(n4342)
         );
  inv0d0 U3485 ( .I(csrbank6_oe0_w[11]), .ZN(n2158) );
  oai22d1 U3486 ( .A1(n2158), .A2(n2181), .B1(n4787), .B2(n2166), .ZN(n4341)
         );
  inv0d0 U3487 ( .I(csrbank6_oe0_w[12]), .ZN(n2159) );
  oai22d1 U3488 ( .A1(n2159), .A2(n2178), .B1(n4598), .B2(n2166), .ZN(n4340)
         );
  inv0d0 U3489 ( .I(csrbank6_oe0_w[13]), .ZN(n2160) );
  oai22d1 U3490 ( .A1(n2160), .A2(n2181), .B1(n5024), .B2(n2180), .ZN(n4339)
         );
  inv0d0 U3491 ( .I(csrbank6_oe0_w[14]), .ZN(n2161) );
  oai22d1 U3492 ( .A1(n2161), .A2(n2181), .B1(n4601), .B2(n2166), .ZN(n4338)
         );
  inv0d0 U3493 ( .I(csrbank6_oe0_w[15]), .ZN(n2162) );
  oai22d1 U3494 ( .A1(n2162), .A2(n2181), .B1(n5028), .B2(n2166), .ZN(n4337)
         );
  inv0d0 U3495 ( .I(csrbank6_oe0_w[16]), .ZN(n2163) );
  oai22d1 U3496 ( .A1(n2163), .A2(n2181), .B1(n2003), .B2(n2166), .ZN(n4336)
         );
  inv0d0 U3497 ( .I(csrbank6_oe0_w[17]), .ZN(n2164) );
  oai22d1 U3498 ( .A1(n2164), .A2(n2178), .B1(n5259), .B2(n2166), .ZN(n4335)
         );
  inv0d0 U3499 ( .I(csrbank6_oe0_w[18]), .ZN(n2165) );
  oai22d1 U3500 ( .A1(n2165), .A2(n2178), .B1(n5260), .B2(n2166), .ZN(n4334)
         );
  inv0d0 U3501 ( .I(csrbank6_oe0_w[19]), .ZN(n2167) );
  oai22d1 U3502 ( .A1(n2167), .A2(n2181), .B1(n5262), .B2(n2166), .ZN(n4333)
         );
  inv0d0 U3503 ( .I(csrbank6_oe0_w[20]), .ZN(n2168) );
  oai22d1 U3504 ( .A1(n2168), .A2(n2181), .B1(n5263), .B2(n2180), .ZN(n4332)
         );
  inv0d0 U3505 ( .I(csrbank6_oe0_w[21]), .ZN(n2169) );
  oai22d1 U3506 ( .A1(n2169), .A2(n2178), .B1(n5264), .B2(n2180), .ZN(n4331)
         );
  inv0d0 U3507 ( .I(csrbank6_oe0_w[22]), .ZN(n2170) );
  oai22d1 U3508 ( .A1(n2170), .A2(n2178), .B1(n5266), .B2(n2180), .ZN(n4330)
         );
  inv0d0 U3509 ( .I(csrbank6_oe0_w[23]), .ZN(n2171) );
  oai22d1 U3510 ( .A1(n2171), .A2(n2178), .B1(n5268), .B2(n2180), .ZN(n4329)
         );
  inv0d0 U3511 ( .I(csrbank6_oe0_w[24]), .ZN(n2172) );
  oai22d1 U3512 ( .A1(n2172), .A2(n2181), .B1(n5270), .B2(n2180), .ZN(n4328)
         );
  inv0d0 U3513 ( .I(csrbank6_oe0_w[25]), .ZN(n2173) );
  oai22d1 U3514 ( .A1(n2173), .A2(n2178), .B1(n5271), .B2(n2180), .ZN(n4327)
         );
  inv0d0 U3515 ( .I(csrbank6_oe0_w[26]), .ZN(n2174) );
  oai22d1 U3516 ( .A1(n2174), .A2(n2181), .B1(n5273), .B2(n2180), .ZN(n4326)
         );
  inv0d0 U3517 ( .I(csrbank6_oe0_w[27]), .ZN(n2175) );
  oai22d1 U3518 ( .A1(n2175), .A2(n2181), .B1(n5275), .B2(n2180), .ZN(n4325)
         );
  inv0d0 U3519 ( .I(csrbank6_oe0_w[28]), .ZN(n2176) );
  oai22d1 U3520 ( .A1(n2176), .A2(n2181), .B1(n5276), .B2(n2180), .ZN(n4324)
         );
  inv0d0 U3521 ( .I(csrbank6_oe0_w[29]), .ZN(n2177) );
  oai22d1 U3522 ( .A1(n2177), .A2(n2178), .B1(n5280), .B2(n2180), .ZN(n4323)
         );
  inv0d0 U3523 ( .I(csrbank6_oe0_w[30]), .ZN(n2179) );
  oai22d1 U3524 ( .A1(n2179), .A2(n2178), .B1(n5283), .B2(n2180), .ZN(n4322)
         );
  inv0d0 U3525 ( .I(csrbank6_oe0_w[31]), .ZN(n2182) );
  oai22d1 U3526 ( .A1(n2182), .A2(n2181), .B1(n5287), .B2(n2180), .ZN(n4321)
         );
  inv0d0 U3527 ( .I(csrbank6_oe1_w[0]), .ZN(n2184) );
  nd02d1 U3528 ( .A1(n5288), .A2(n2186), .ZN(n2210) );
  aoi22d1 U3529 ( .A1(n2184), .A2(n2186), .B1(n5000), .B2(n2210), .ZN(n4320)
         );
  inv0d0 U3530 ( .I(csrbank6_oe1_w[1]), .ZN(n2185) );
  aoi22d1 U3531 ( .A1(n2185), .A2(n2186), .B1(n2653), .B2(n2210), .ZN(n4319)
         );
  inv0d0 U3532 ( .I(csrbank6_oe1_w[2]), .ZN(n2187) );
  or02d1 U3533 ( .A1(n2186), .A2(n5111), .Z(n2216) );
  buffd1 U3534 ( .I(n2216), .Z(n2218) );
  oai22d1 U3535 ( .A1(n2187), .A2(n2210), .B1(n5004), .B2(n2218), .ZN(n4318)
         );
  inv0d0 U3536 ( .I(csrbank6_oe1_w[3]), .ZN(n2188) );
  oai22d1 U3537 ( .A1(n2188), .A2(n2210), .B1(n5246), .B2(n2218), .ZN(n4317)
         );
  inv0d0 U3538 ( .I(csrbank6_oe1_w[4]), .ZN(n2189) );
  buffd1 U3539 ( .I(n2210), .Z(n2219) );
  oai22d1 U3540 ( .A1(n2189), .A2(n2219), .B1(n5247), .B2(n2218), .ZN(n4316)
         );
  inv0d0 U3541 ( .I(csrbank6_oe1_w[5]), .ZN(n2190) );
  oai22d1 U3542 ( .A1(n2190), .A2(n2210), .B1(n5248), .B2(n2218), .ZN(n4315)
         );
  inv0d0 U3543 ( .I(csrbank6_oe1_w[6]), .ZN(n2191) );
  oai22d1 U3544 ( .A1(n2191), .A2(n2210), .B1(n5249), .B2(n2218), .ZN(n4314)
         );
  inv0d0 U3545 ( .I(csrbank6_oe1_w[7]), .ZN(n2192) );
  oai22d1 U3546 ( .A1(n2192), .A2(n2210), .B1(n2635), .B2(n2218), .ZN(n4313)
         );
  inv0d0 U3547 ( .I(csrbank6_oe1_w[8]), .ZN(n2193) );
  oai22d1 U3548 ( .A1(n2193), .A2(n2219), .B1(n4783), .B2(n2218), .ZN(n4312)
         );
  inv0d0 U3549 ( .I(csrbank6_oe1_w[9]), .ZN(n2194) );
  oai22d1 U3550 ( .A1(n2194), .A2(n2219), .B1(n4593), .B2(n2218), .ZN(n4311)
         );
  inv0d0 U3551 ( .I(csrbank6_oe1_w[10]), .ZN(n2195) );
  oai22d1 U3552 ( .A1(n2195), .A2(n2210), .B1(n4595), .B2(n2218), .ZN(n4310)
         );
  inv0d0 U3553 ( .I(csrbank6_oe1_w[11]), .ZN(n2196) );
  oai22d1 U3554 ( .A1(n2196), .A2(n2210), .B1(n5254), .B2(n2216), .ZN(n4309)
         );
  inv0d0 U3555 ( .I(csrbank6_oe1_w[12]), .ZN(n2197) );
  oai22d1 U3556 ( .A1(n2197), .A2(n2219), .B1(n4598), .B2(n2216), .ZN(n4308)
         );
  inv0d0 U3557 ( .I(csrbank6_oe1_w[13]), .ZN(n2198) );
  oai22d1 U3558 ( .A1(n2198), .A2(n2210), .B1(n4790), .B2(n2216), .ZN(n4307)
         );
  inv0d0 U3559 ( .I(csrbank6_oe1_w[14]), .ZN(n2199) );
  oai22d1 U3560 ( .A1(n2199), .A2(n2210), .B1(n4601), .B2(n2216), .ZN(n4306)
         );
  inv0d0 U3561 ( .I(csrbank6_oe1_w[15]), .ZN(n2200) );
  oai22d1 U3562 ( .A1(n2200), .A2(n2210), .B1(n4793), .B2(n2216), .ZN(n4305)
         );
  inv0d0 U3563 ( .I(csrbank6_oe1_w[16]), .ZN(n2201) );
  oai22d1 U3564 ( .A1(n2201), .A2(n2219), .B1(n2003), .B2(n2216), .ZN(n4304)
         );
  inv0d0 U3565 ( .I(csrbank6_oe1_w[17]), .ZN(n2202) );
  oai22d1 U3566 ( .A1(n2202), .A2(n2219), .B1(n5259), .B2(n2216), .ZN(n4303)
         );
  inv0d0 U3567 ( .I(csrbank6_oe1_w[18]), .ZN(n2203) );
  oai22d1 U3568 ( .A1(n2203), .A2(n2219), .B1(n5260), .B2(n2218), .ZN(n4302)
         );
  inv0d0 U3569 ( .I(csrbank6_oe1_w[19]), .ZN(n2204) );
  oai22d1 U3570 ( .A1(n2204), .A2(n2219), .B1(n5262), .B2(n2216), .ZN(n4301)
         );
  inv0d0 U3571 ( .I(csrbank6_oe1_w[20]), .ZN(n2205) );
  oai22d1 U3572 ( .A1(n2205), .A2(n2219), .B1(n5263), .B2(n2216), .ZN(n4300)
         );
  inv0d0 U3573 ( .I(csrbank6_oe1_w[21]), .ZN(n2206) );
  oai22d1 U3574 ( .A1(n2206), .A2(n2219), .B1(n5264), .B2(n2216), .ZN(n4299)
         );
  inv0d0 U3575 ( .I(csrbank6_oe1_w[22]), .ZN(n2207) );
  oai22d1 U3576 ( .A1(n2207), .A2(n2210), .B1(n5266), .B2(n2216), .ZN(n4298)
         );
  inv0d0 U3577 ( .I(csrbank6_oe1_w[23]), .ZN(n2208) );
  oai22d1 U3578 ( .A1(n2208), .A2(n2219), .B1(n5268), .B2(n2218), .ZN(n4297)
         );
  inv0d0 U3579 ( .I(csrbank6_oe1_w[24]), .ZN(n2209) );
  oai22d1 U3580 ( .A1(n2209), .A2(n2210), .B1(n5270), .B2(n2218), .ZN(n4296)
         );
  inv0d0 U3581 ( .I(csrbank6_oe1_w[25]), .ZN(n2211) );
  oai22d1 U3582 ( .A1(n2211), .A2(n2210), .B1(n5271), .B2(n2218), .ZN(n4295)
         );
  inv0d0 U3583 ( .I(csrbank6_oe1_w[26]), .ZN(n2212) );
  oai22d1 U3584 ( .A1(n2212), .A2(n2219), .B1(n5273), .B2(n2218), .ZN(n4294)
         );
  inv0d0 U3585 ( .I(csrbank6_oe1_w[27]), .ZN(n2213) );
  oai22d1 U3586 ( .A1(n2213), .A2(n2219), .B1(n5275), .B2(n2218), .ZN(n4293)
         );
  inv0d0 U3587 ( .I(csrbank6_oe1_w[28]), .ZN(n2214) );
  oai22d1 U3588 ( .A1(n2214), .A2(n2219), .B1(n5276), .B2(n2216), .ZN(n4292)
         );
  inv0d0 U3589 ( .I(csrbank6_oe1_w[29]), .ZN(n2215) );
  oai22d1 U3590 ( .A1(n2215), .A2(n2219), .B1(n5280), .B2(n2218), .ZN(n4291)
         );
  inv0d0 U3591 ( .I(csrbank6_oe1_w[30]), .ZN(n2217) );
  oai22d1 U3592 ( .A1(n2217), .A2(n2219), .B1(n5283), .B2(n2216), .ZN(n4290)
         );
  inv0d0 U3593 ( .I(csrbank6_oe1_w[31]), .ZN(n2220) );
  oai22d1 U3594 ( .A1(n2220), .A2(n2219), .B1(n5287), .B2(n2218), .ZN(n4289)
         );
  inv0d0 U3595 ( .I(csrbank6_oe2_w[0]), .ZN(n2222) );
  oaim21d1 U3596 ( .B1(n4683), .B2(n2221), .A(n5956), .ZN(n2248) );
  nd02d1 U3597 ( .A1(n2221), .A2(n4580), .ZN(n2255) );
  buffd1 U3598 ( .I(n2255), .Z(n2253) );
  oai22d1 U3599 ( .A1(n2222), .A2(n2248), .B1(n5290), .B2(n2253), .ZN(n4288)
         );
  inv0d0 U3600 ( .I(csrbank6_oe2_w[1]), .ZN(n2223) );
  oai22d1 U3601 ( .A1(n2223), .A2(n2248), .B1(n2639), .B2(n2253), .ZN(n4287)
         );
  inv0d0 U3602 ( .I(csrbank6_oe2_w[2]), .ZN(n2224) );
  oai22d1 U3603 ( .A1(n2224), .A2(n2248), .B1(n5004), .B2(n2253), .ZN(n4286)
         );
  inv0d0 U3604 ( .I(csrbank6_oe2_w[3]), .ZN(n2225) );
  oai22d1 U3605 ( .A1(n2225), .A2(n2248), .B1(n5246), .B2(n2253), .ZN(n4285)
         );
  inv0d0 U3606 ( .I(csrbank6_oe2_w[4]), .ZN(n2226) );
  buffd1 U3607 ( .I(n2248), .Z(n2256) );
  oai22d1 U3608 ( .A1(n2226), .A2(n2256), .B1(n5247), .B2(n2253), .ZN(n4284)
         );
  inv0d0 U3609 ( .I(csrbank6_oe2_w[5]), .ZN(n2227) );
  oai22d1 U3610 ( .A1(n2227), .A2(n2248), .B1(n5248), .B2(n2253), .ZN(n4283)
         );
  inv0d0 U3611 ( .I(csrbank6_oe2_w[6]), .ZN(n2228) );
  oai22d1 U3612 ( .A1(n2228), .A2(n2248), .B1(n5249), .B2(n2253), .ZN(n4282)
         );
  inv0d0 U3613 ( .I(csrbank6_oe2_w[7]), .ZN(n2229) );
  oai22d1 U3614 ( .A1(n2229), .A2(n2248), .B1(n2635), .B2(n2253), .ZN(n4281)
         );
  inv0d0 U3615 ( .I(csrbank6_oe2_w[8]), .ZN(n2230) );
  oai22d1 U3616 ( .A1(n2230), .A2(n2248), .B1(n4783), .B2(n2253), .ZN(n4280)
         );
  inv0d0 U3617 ( .I(csrbank6_oe2_w[9]), .ZN(n2231) );
  oai22d1 U3618 ( .A1(n2231), .A2(n2256), .B1(n4593), .B2(n2253), .ZN(n4279)
         );
  inv0d0 U3619 ( .I(csrbank6_oe2_w[10]), .ZN(n2232) );
  oai22d1 U3620 ( .A1(n2232), .A2(n2256), .B1(n4595), .B2(n2255), .ZN(n4278)
         );
  inv0d0 U3621 ( .I(csrbank6_oe2_w[11]), .ZN(n2233) );
  oai22d1 U3622 ( .A1(n2233), .A2(n2256), .B1(n5254), .B2(n2255), .ZN(n4277)
         );
  inv0d0 U3623 ( .I(csrbank6_oe2_w[12]), .ZN(n2234) );
  oai22d1 U3624 ( .A1(n2234), .A2(n2256), .B1(n4598), .B2(n2255), .ZN(n4276)
         );
  inv0d0 U3625 ( .I(csrbank6_oe2_w[13]), .ZN(n2235) );
  oai22d1 U3626 ( .A1(n2235), .A2(n2256), .B1(n4790), .B2(n2253), .ZN(n4275)
         );
  inv0d0 U3627 ( .I(csrbank6_oe2_w[14]), .ZN(n2236) );
  oai22d1 U3628 ( .A1(n2236), .A2(n2256), .B1(n4601), .B2(n2253), .ZN(n4274)
         );
  inv0d0 U3629 ( .I(csrbank6_oe2_w[15]), .ZN(n2237) );
  oai22d1 U3630 ( .A1(n2237), .A2(n2256), .B1(n4793), .B2(n2255), .ZN(n4273)
         );
  inv0d0 U3631 ( .I(csrbank6_oe2_w[16]), .ZN(n2238) );
  oai22d1 U3632 ( .A1(n2238), .A2(n2248), .B1(n2003), .B2(n2255), .ZN(n4272)
         );
  inv0d0 U3633 ( .I(csrbank6_oe2_w[17]), .ZN(n2239) );
  oai22d1 U3634 ( .A1(n2239), .A2(n2248), .B1(n5259), .B2(n2253), .ZN(n4271)
         );
  inv0d0 U3635 ( .I(csrbank6_oe2_w[18]), .ZN(n2240) );
  oai22d1 U3636 ( .A1(n2240), .A2(n2256), .B1(n5260), .B2(n2255), .ZN(n4270)
         );
  inv0d0 U3637 ( .I(csrbank6_oe2_w[19]), .ZN(n2241) );
  oai22d1 U3638 ( .A1(n2241), .A2(n2248), .B1(n5262), .B2(n2255), .ZN(n4269)
         );
  inv0d0 U3639 ( .I(csrbank6_oe2_w[20]), .ZN(n2242) );
  oai22d1 U3640 ( .A1(n2242), .A2(n2248), .B1(n5263), .B2(n2255), .ZN(n4268)
         );
  inv0d0 U3641 ( .I(csrbank6_oe2_w[21]), .ZN(n2243) );
  oai22d1 U3642 ( .A1(n2243), .A2(n2248), .B1(n5264), .B2(n2255), .ZN(n4267)
         );
  inv0d0 U3643 ( .I(csrbank6_oe2_w[22]), .ZN(n2244) );
  oai22d1 U3644 ( .A1(n2244), .A2(n2248), .B1(n5266), .B2(n2255), .ZN(n4266)
         );
  inv0d0 U3645 ( .I(csrbank6_oe2_w[23]), .ZN(n2245) );
  oai22d1 U3646 ( .A1(n2245), .A2(n2248), .B1(n5268), .B2(n2255), .ZN(n4265)
         );
  inv0d0 U3647 ( .I(csrbank6_oe2_w[24]), .ZN(n2246) );
  oai22d1 U3648 ( .A1(n2246), .A2(n2256), .B1(n5270), .B2(n2255), .ZN(n4264)
         );
  inv0d0 U3649 ( .I(csrbank6_oe2_w[25]), .ZN(n2247) );
  oai22d1 U3650 ( .A1(n2247), .A2(n2256), .B1(n5271), .B2(n2255), .ZN(n4263)
         );
  inv0d0 U3651 ( .I(csrbank6_oe2_w[26]), .ZN(n2249) );
  oai22d1 U3652 ( .A1(n2249), .A2(n2248), .B1(n5273), .B2(n2255), .ZN(n4262)
         );
  inv0d0 U3653 ( .I(csrbank6_oe2_w[27]), .ZN(n2250) );
  oai22d1 U3654 ( .A1(n2250), .A2(n2256), .B1(n5275), .B2(n2253), .ZN(n4261)
         );
  inv0d0 U3655 ( .I(csrbank6_oe2_w[28]), .ZN(n2251) );
  oai22d1 U3656 ( .A1(n2251), .A2(n2256), .B1(n5276), .B2(n2253), .ZN(n4260)
         );
  inv0d0 U3657 ( .I(csrbank6_oe2_w[29]), .ZN(n2252) );
  oai22d1 U3658 ( .A1(n2252), .A2(n2256), .B1(n5280), .B2(n2253), .ZN(n4259)
         );
  inv0d0 U3659 ( .I(csrbank6_oe2_w[30]), .ZN(n2254) );
  oai22d1 U3660 ( .A1(n2254), .A2(n2256), .B1(n5283), .B2(n2253), .ZN(n4258)
         );
  inv0d0 U3661 ( .I(csrbank6_oe2_w[31]), .ZN(n2257) );
  oai22d1 U3662 ( .A1(n2257), .A2(n2256), .B1(n5287), .B2(n2255), .ZN(n4257)
         );
  inv0d0 U3663 ( .I(csrbank6_oe3_w[0]), .ZN(n2259) );
  oai21d1 U3664 ( .B1(n2372), .B2(n2654), .A(n5319), .ZN(n2285) );
  nd03d1 U3665 ( .A1(n2373), .A2(n2258), .A3(n5301), .ZN(n2292) );
  buffd1 U3666 ( .I(n2292), .Z(n2290) );
  oai22d1 U3667 ( .A1(n2259), .A2(n2285), .B1(n266), .B2(n2290), .ZN(n4256) );
  inv0d0 U3668 ( .I(csrbank6_oe3_w[1]), .ZN(n2260) );
  oai22d1 U3669 ( .A1(n2260), .A2(n2285), .B1(n2639), .B2(n2290), .ZN(n4255)
         );
  inv0d0 U3670 ( .I(csrbank6_oe3_w[2]), .ZN(n2261) );
  oai22d1 U3671 ( .A1(n2261), .A2(n2285), .B1(n5004), .B2(n2290), .ZN(n4254)
         );
  inv0d0 U3672 ( .I(csrbank6_oe3_w[3]), .ZN(n2262) );
  oai22d1 U3673 ( .A1(n2262), .A2(n2285), .B1(n5246), .B2(n2290), .ZN(n4253)
         );
  inv0d0 U3674 ( .I(csrbank6_oe3_w[4]), .ZN(n2263) );
  buffd1 U3675 ( .I(n2285), .Z(n2293) );
  oai22d1 U3676 ( .A1(n2263), .A2(n2293), .B1(n5247), .B2(n2290), .ZN(n4252)
         );
  inv0d0 U3677 ( .I(csrbank6_oe3_w[5]), .ZN(n2264) );
  oai22d1 U3678 ( .A1(n2264), .A2(n2293), .B1(n5248), .B2(n2290), .ZN(n4251)
         );
  inv0d0 U3679 ( .I(csrbank6_oe3_w[6]), .ZN(n2265) );
  oai22d1 U3680 ( .A1(n2265), .A2(n2285), .B1(n5249), .B2(n2290), .ZN(n4250)
         );
  inv0d0 U3681 ( .I(csrbank6_oe3_w[7]), .ZN(n2266) );
  oai22d1 U3682 ( .A1(n2266), .A2(n2285), .B1(n2635), .B2(n2290), .ZN(n4249)
         );
  inv0d0 U3683 ( .I(csrbank6_oe3_w[8]), .ZN(n2267) );
  oai22d1 U3684 ( .A1(n2267), .A2(n2285), .B1(n4783), .B2(n2290), .ZN(n4248)
         );
  inv0d0 U3685 ( .I(csrbank6_oe3_w[9]), .ZN(n2268) );
  oai22d1 U3686 ( .A1(n2268), .A2(n2293), .B1(n4593), .B2(n2292), .ZN(n4247)
         );
  inv0d0 U3687 ( .I(csrbank6_oe3_w[10]), .ZN(n2269) );
  oai22d1 U3688 ( .A1(n2269), .A2(n2285), .B1(n4595), .B2(n2290), .ZN(n4246)
         );
  inv0d0 U3689 ( .I(csrbank6_oe3_w[11]), .ZN(n2270) );
  oai22d1 U3690 ( .A1(n2270), .A2(n2285), .B1(n5254), .B2(n2290), .ZN(n4245)
         );
  inv0d0 U3691 ( .I(csrbank6_oe3_w[12]), .ZN(n2271) );
  oai22d1 U3692 ( .A1(n2271), .A2(n2293), .B1(n4598), .B2(n2290), .ZN(n4244)
         );
  inv0d0 U3693 ( .I(csrbank6_oe3_w[13]), .ZN(n2272) );
  oai22d1 U3694 ( .A1(n2272), .A2(n2285), .B1(n4790), .B2(n2292), .ZN(n4243)
         );
  inv0d0 U3695 ( .I(csrbank6_oe3_w[14]), .ZN(n2273) );
  oai22d1 U3696 ( .A1(n2273), .A2(n2285), .B1(n4601), .B2(n2292), .ZN(n4242)
         );
  inv0d0 U3697 ( .I(csrbank6_oe3_w[15]), .ZN(n2274) );
  oai22d1 U3698 ( .A1(n2274), .A2(n2293), .B1(n4793), .B2(n2292), .ZN(n4241)
         );
  inv0d0 U3699 ( .I(csrbank6_oe3_w[16]), .ZN(n2275) );
  oai22d1 U3700 ( .A1(n2275), .A2(n2293), .B1(n2003), .B2(n2290), .ZN(n4240)
         );
  inv0d0 U3701 ( .I(csrbank6_oe3_w[17]), .ZN(n2276) );
  oai22d1 U3702 ( .A1(n2276), .A2(n2293), .B1(n5259), .B2(n2292), .ZN(n4239)
         );
  inv0d0 U3703 ( .I(csrbank6_oe3_w[18]), .ZN(n2277) );
  oai22d1 U3704 ( .A1(n2277), .A2(n2293), .B1(n5260), .B2(n2292), .ZN(n4238)
         );
  inv0d0 U3705 ( .I(csrbank6_oe3_w[19]), .ZN(n2278) );
  oai22d1 U3706 ( .A1(n2278), .A2(n2293), .B1(n5262), .B2(n2292), .ZN(n4237)
         );
  inv0d0 U3707 ( .I(csrbank6_oe3_w[20]), .ZN(n2279) );
  oai22d1 U3708 ( .A1(n2279), .A2(n2285), .B1(n5263), .B2(n2292), .ZN(n4236)
         );
  inv0d0 U3709 ( .I(csrbank6_oe3_w[21]), .ZN(n2280) );
  oai22d1 U3710 ( .A1(n2280), .A2(n2293), .B1(n5264), .B2(n2292), .ZN(n4235)
         );
  inv0d0 U3711 ( .I(csrbank6_oe3_w[22]), .ZN(n2281) );
  oai22d1 U3712 ( .A1(n2281), .A2(n2285), .B1(n5266), .B2(n2292), .ZN(n4234)
         );
  inv0d0 U3713 ( .I(csrbank6_oe3_w[23]), .ZN(n2282) );
  oai22d1 U3714 ( .A1(n2282), .A2(n2293), .B1(n5268), .B2(n2292), .ZN(n4233)
         );
  inv0d0 U3715 ( .I(csrbank6_oe3_w[24]), .ZN(n2283) );
  oai22d1 U3716 ( .A1(n2283), .A2(n2293), .B1(n5270), .B2(n2292), .ZN(n4232)
         );
  inv0d0 U3717 ( .I(csrbank6_oe3_w[25]), .ZN(n2284) );
  oai22d1 U3718 ( .A1(n2284), .A2(n2285), .B1(n5271), .B2(n2292), .ZN(n4231)
         );
  inv0d0 U3719 ( .I(csrbank6_oe3_w[26]), .ZN(n2286) );
  oai22d1 U3720 ( .A1(n2286), .A2(n2285), .B1(n5273), .B2(n2292), .ZN(n4230)
         );
  inv0d0 U3721 ( .I(csrbank6_oe3_w[27]), .ZN(n2287) );
  oai22d1 U3722 ( .A1(n2287), .A2(n2293), .B1(n5275), .B2(n2290), .ZN(n4229)
         );
  inv0d0 U3723 ( .I(csrbank6_oe3_w[28]), .ZN(n2288) );
  oai22d1 U3724 ( .A1(n2288), .A2(n2293), .B1(n5276), .B2(n2290), .ZN(n4228)
         );
  inv0d0 U3725 ( .I(csrbank6_oe3_w[29]), .ZN(n2289) );
  oai22d1 U3726 ( .A1(n2289), .A2(n2293), .B1(n5280), .B2(n2290), .ZN(n4227)
         );
  inv0d0 U3727 ( .I(csrbank6_oe3_w[30]), .ZN(n2291) );
  oai22d1 U3728 ( .A1(n2291), .A2(n2293), .B1(n5283), .B2(n2290), .ZN(n4226)
         );
  inv0d0 U3729 ( .I(csrbank6_oe3_w[31]), .ZN(n2294) );
  oai22d1 U3730 ( .A1(n2294), .A2(n2293), .B1(n5287), .B2(n2292), .ZN(n4225)
         );
  inv0d0 U3731 ( .I(csrbank6_ien0_w[0]), .ZN(n2296) );
  nd02d1 U3732 ( .A1(n5288), .A2(n2300), .ZN(n2323) );
  aoi22d1 U3733 ( .A1(n2296), .A2(n2300), .B1(n4955), .B2(n2323), .ZN(n4224)
         );
  inv0d0 U3734 ( .I(csrbank6_ien0_w[1]), .ZN(n2297) );
  aoi22d1 U3735 ( .A1(n2297), .A2(n2300), .B1(n2653), .B2(n2323), .ZN(n4223)
         );
  inv0d0 U3736 ( .I(csrbank6_ien0_w[2]), .ZN(n2299) );
  aoi22d1 U3737 ( .A1(n2299), .A2(n2300), .B1(n2298), .B2(n2323), .ZN(n4222)
         );
  inv0d0 U3738 ( .I(csrbank6_ien0_w[3]), .ZN(n2301) );
  oai22d1 U3739 ( .A1(n2301), .A2(n2323), .B1(n5246), .B2(n2328), .ZN(n4221)
         );
  inv0d0 U3740 ( .I(csrbank6_ien0_w[4]), .ZN(n2302) );
  buffd1 U3741 ( .I(n2323), .Z(n2332) );
  oai22d1 U3742 ( .A1(n2302), .A2(n2332), .B1(n5247), .B2(n2328), .ZN(n4220)
         );
  inv0d0 U3743 ( .I(csrbank6_ien0_w[5]), .ZN(n2303) );
  oai22d1 U3744 ( .A1(n2303), .A2(n2323), .B1(n5248), .B2(n2328), .ZN(n4219)
         );
  inv0d0 U3745 ( .I(csrbank6_ien0_w[6]), .ZN(n2304) );
  oai22d1 U3746 ( .A1(n2304), .A2(n2323), .B1(n5012), .B2(n2328), .ZN(n4218)
         );
  inv0d0 U3747 ( .I(csrbank6_ien0_w[7]), .ZN(n2305) );
  oai22d1 U3748 ( .A1(n2305), .A2(n2323), .B1(n5251), .B2(n2328), .ZN(n4217)
         );
  inv0d0 U3749 ( .I(csrbank6_ien0_w[8]), .ZN(n2306) );
  oai22d1 U3750 ( .A1(n2306), .A2(n2323), .B1(n5015), .B2(n2328), .ZN(n4216)
         );
  inv0d0 U3751 ( .I(csrbank6_ien0_w[9]), .ZN(n2307) );
  oai22d1 U3752 ( .A1(n2307), .A2(n2332), .B1(n5017), .B2(n2328), .ZN(n4215)
         );
  inv0d0 U3753 ( .I(csrbank6_ien0_w[10]), .ZN(n2308) );
  oai22d1 U3754 ( .A1(n2308), .A2(n2323), .B1(n5019), .B2(n2328), .ZN(n4214)
         );
  inv0d0 U3755 ( .I(csrbank6_ien0_w[11]), .ZN(n2309) );
  oai22d1 U3756 ( .A1(n2309), .A2(n2323), .B1(n4787), .B2(n2328), .ZN(n4213)
         );
  inv0d0 U3757 ( .I(csrbank6_ien0_w[12]), .ZN(n2310) );
  oai22d1 U3758 ( .A1(n2310), .A2(n2332), .B1(n5022), .B2(n2328), .ZN(n4212)
         );
  inv0d0 U3759 ( .I(csrbank6_ien0_w[13]), .ZN(n2311) );
  oai22d1 U3760 ( .A1(n2311), .A2(n2323), .B1(n5024), .B2(n2328), .ZN(n4211)
         );
  inv0d0 U3761 ( .I(csrbank6_ien0_w[14]), .ZN(n2312) );
  oai22d1 U3762 ( .A1(n2312), .A2(n2323), .B1(n5026), .B2(n2328), .ZN(n4210)
         );
  inv0d0 U3763 ( .I(csrbank6_ien0_w[15]), .ZN(n2313) );
  oai22d1 U3764 ( .A1(n2313), .A2(n2332), .B1(n5028), .B2(n2328), .ZN(n4209)
         );
  inv0d0 U3765 ( .I(csrbank6_ien0_w[16]), .ZN(n2314) );
  oai22d1 U3766 ( .A1(n2314), .A2(n2332), .B1(n2003), .B2(n2328), .ZN(n4208)
         );
  inv0d0 U3767 ( .I(csrbank6_ien0_w[17]), .ZN(n2315) );
  oai22d1 U3768 ( .A1(n2315), .A2(n2332), .B1(n5259), .B2(n2328), .ZN(n4207)
         );
  inv0d0 U3769 ( .I(csrbank6_ien0_w[18]), .ZN(n2316) );
  oai22d1 U3770 ( .A1(n2316), .A2(n2332), .B1(n5260), .B2(n2328), .ZN(n4206)
         );
  inv0d0 U3771 ( .I(csrbank6_ien0_w[19]), .ZN(n2317) );
  oai22d1 U3772 ( .A1(n2317), .A2(n2332), .B1(n5262), .B2(n2328), .ZN(n4205)
         );
  inv0d0 U3773 ( .I(csrbank6_ien0_w[20]), .ZN(n2318) );
  oai22d1 U3774 ( .A1(n2318), .A2(n2332), .B1(n5263), .B2(n2328), .ZN(n4204)
         );
  inv0d0 U3775 ( .I(csrbank6_ien0_w[21]), .ZN(n2319) );
  oai22d1 U3776 ( .A1(n2319), .A2(n2332), .B1(n5264), .B2(n2328), .ZN(n4203)
         );
  inv0d0 U3777 ( .I(csrbank6_ien0_w[22]), .ZN(n2320) );
  oai22d1 U3778 ( .A1(n2320), .A2(n2323), .B1(n5266), .B2(n2328), .ZN(n4202)
         );
  inv0d0 U3779 ( .I(csrbank6_ien0_w[23]), .ZN(n2321) );
  oai22d1 U3780 ( .A1(n2321), .A2(n2332), .B1(n5268), .B2(n2328), .ZN(n4201)
         );
  inv0d0 U3781 ( .I(csrbank6_ien0_w[24]), .ZN(n2322) );
  oai22d1 U3782 ( .A1(n2322), .A2(n2323), .B1(n5270), .B2(n2328), .ZN(n4200)
         );
  inv0d0 U3783 ( .I(csrbank6_ien0_w[25]), .ZN(n2324) );
  oai22d1 U3784 ( .A1(n2324), .A2(n2323), .B1(n5271), .B2(n2328), .ZN(n4199)
         );
  inv0d0 U3785 ( .I(csrbank6_ien0_w[26]), .ZN(n2325) );
  oai22d1 U3786 ( .A1(n2325), .A2(n2332), .B1(n5273), .B2(n2328), .ZN(n4198)
         );
  inv0d0 U3787 ( .I(csrbank6_ien0_w[27]), .ZN(n2326) );
  oai22d1 U3788 ( .A1(n2326), .A2(n2332), .B1(n5275), .B2(n2328), .ZN(n4197)
         );
  inv0d0 U3789 ( .I(csrbank6_ien0_w[28]), .ZN(n2327) );
  oai22d1 U3790 ( .A1(n2327), .A2(n2332), .B1(n5276), .B2(n2328), .ZN(n4196)
         );
  inv0d0 U3791 ( .I(csrbank6_ien0_w[29]), .ZN(n2329) );
  oai22d1 U3792 ( .A1(n2329), .A2(n2332), .B1(n5280), .B2(n2328), .ZN(n4195)
         );
  inv0d0 U3793 ( .I(csrbank6_ien0_w[30]), .ZN(n2330) );
  oai22d1 U3794 ( .A1(n2330), .A2(n2332), .B1(n5283), .B2(n2328), .ZN(n4194)
         );
  inv0d0 U3795 ( .I(csrbank6_ien0_w[31]), .ZN(n2333) );
  oai22d1 U3796 ( .A1(n2333), .A2(n2332), .B1(n5287), .B2(n2328), .ZN(n4193)
         );
  inv0d0 U3797 ( .I(csrbank6_ien1_w[0]), .ZN(n2336) );
  oai21d1 U3798 ( .B1(n2372), .B2(n2334), .A(n5955), .ZN(n2362) );
  nd03d1 U3799 ( .A1(n2373), .A2(n2335), .A3(n5288), .ZN(n2369) );
  buffd1 U3800 ( .I(n2369), .Z(n2367) );
  oai22d1 U3801 ( .A1(n2336), .A2(n2362), .B1(n4808), .B2(n2367), .ZN(n4192)
         );
  inv0d0 U3802 ( .I(csrbank6_ien1_w[1]), .ZN(n2337) );
  oai22d1 U3803 ( .A1(n2337), .A2(n2362), .B1(n2639), .B2(n2367), .ZN(n4191)
         );
  inv0d0 U3804 ( .I(csrbank6_ien1_w[2]), .ZN(n2338) );
  oai22d1 U3805 ( .A1(n2338), .A2(n2362), .B1(n5004), .B2(n2367), .ZN(n4190)
         );
  inv0d0 U3806 ( .I(csrbank6_ien1_w[3]), .ZN(n2339) );
  oai22d1 U3807 ( .A1(n2339), .A2(n2362), .B1(n2625), .B2(n2367), .ZN(n4189)
         );
  inv0d0 U3808 ( .I(csrbank6_ien1_w[4]), .ZN(n2340) );
  buffd1 U3809 ( .I(n2362), .Z(n2370) );
  oai22d1 U3810 ( .A1(n2340), .A2(n2370), .B1(n5247), .B2(n2367), .ZN(n4188)
         );
  inv0d0 U3811 ( .I(csrbank6_ien1_w[5]), .ZN(n2341) );
  oai22d1 U3812 ( .A1(n2341), .A2(n2370), .B1(n5010), .B2(n2367), .ZN(n4187)
         );
  inv0d0 U3813 ( .I(csrbank6_ien1_w[6]), .ZN(n2342) );
  oai22d1 U3814 ( .A1(n2342), .A2(n2362), .B1(n5012), .B2(n2367), .ZN(n4186)
         );
  inv0d0 U3815 ( .I(csrbank6_ien1_w[7]), .ZN(n2343) );
  oai22d1 U3816 ( .A1(n2343), .A2(n2362), .B1(n2635), .B2(n2367), .ZN(n4185)
         );
  inv0d0 U3817 ( .I(csrbank6_ien1_w[8]), .ZN(n2344) );
  oai22d1 U3818 ( .A1(n2344), .A2(n2362), .B1(n5015), .B2(n2367), .ZN(n4184)
         );
  inv0d0 U3819 ( .I(csrbank6_ien1_w[9]), .ZN(n2345) );
  oai22d1 U3820 ( .A1(n2345), .A2(n2370), .B1(n5017), .B2(n2369), .ZN(n4183)
         );
  inv0d0 U3821 ( .I(csrbank6_ien1_w[10]), .ZN(n2346) );
  oai22d1 U3822 ( .A1(n2346), .A2(n2362), .B1(n5019), .B2(n2367), .ZN(n4182)
         );
  inv0d0 U3823 ( .I(csrbank6_ien1_w[11]), .ZN(n2347) );
  oai22d1 U3824 ( .A1(n2347), .A2(n2362), .B1(n4787), .B2(n2367), .ZN(n4181)
         );
  inv0d0 U3825 ( .I(csrbank6_ien1_w[12]), .ZN(n2348) );
  oai22d1 U3826 ( .A1(n2348), .A2(n2370), .B1(n5022), .B2(n2367), .ZN(n4180)
         );
  inv0d0 U3827 ( .I(csrbank6_ien1_w[13]), .ZN(n2349) );
  oai22d1 U3828 ( .A1(n2349), .A2(n2362), .B1(n5024), .B2(n2369), .ZN(n4179)
         );
  inv0d0 U3829 ( .I(csrbank6_ien1_w[14]), .ZN(n2350) );
  oai22d1 U3830 ( .A1(n2350), .A2(n2362), .B1(n5026), .B2(n2369), .ZN(n4178)
         );
  inv0d0 U3831 ( .I(csrbank6_ien1_w[15]), .ZN(n2351) );
  oai22d1 U3832 ( .A1(n2351), .A2(n2370), .B1(n5028), .B2(n2369), .ZN(n4177)
         );
  inv0d0 U3833 ( .I(csrbank6_ien1_w[16]), .ZN(n2352) );
  oai22d1 U3834 ( .A1(n2352), .A2(n2370), .B1(n2003), .B2(n2367), .ZN(n4176)
         );
  inv0d0 U3835 ( .I(csrbank6_ien1_w[17]), .ZN(n2353) );
  oai22d1 U3836 ( .A1(n2353), .A2(n2370), .B1(n5259), .B2(n2369), .ZN(n4175)
         );
  inv0d0 U3837 ( .I(csrbank6_ien1_w[18]), .ZN(n2354) );
  oai22d1 U3838 ( .A1(n2354), .A2(n2362), .B1(n5260), .B2(n2369), .ZN(n4174)
         );
  inv0d0 U3839 ( .I(csrbank6_ien1_w[19]), .ZN(n2355) );
  oai22d1 U3840 ( .A1(n2355), .A2(n2370), .B1(n5262), .B2(n2369), .ZN(n4173)
         );
  inv0d0 U3841 ( .I(csrbank6_ien1_w[20]), .ZN(n2356) );
  oai22d1 U3842 ( .A1(n2356), .A2(n2362), .B1(n5263), .B2(n2369), .ZN(n4172)
         );
  inv0d0 U3843 ( .I(csrbank6_ien1_w[21]), .ZN(n2357) );
  oai22d1 U3844 ( .A1(n2357), .A2(n2370), .B1(n5264), .B2(n2369), .ZN(n4171)
         );
  inv0d0 U3845 ( .I(csrbank6_ien1_w[22]), .ZN(n2358) );
  oai22d1 U3846 ( .A1(n2358), .A2(n2362), .B1(n5266), .B2(n2369), .ZN(n4170)
         );
  inv0d0 U3847 ( .I(csrbank6_ien1_w[23]), .ZN(n2359) );
  oai22d1 U3848 ( .A1(n2359), .A2(n2370), .B1(n5268), .B2(n2369), .ZN(n4169)
         );
  inv0d0 U3849 ( .I(csrbank6_ien1_w[24]), .ZN(n2360) );
  oai22d1 U3850 ( .A1(n2360), .A2(n2370), .B1(n5270), .B2(n2369), .ZN(n4168)
         );
  inv0d0 U3851 ( .I(csrbank6_ien1_w[25]), .ZN(n2361) );
  oai22d1 U3852 ( .A1(n2361), .A2(n2370), .B1(n5271), .B2(n2369), .ZN(n4167)
         );
  inv0d0 U3853 ( .I(csrbank6_ien1_w[26]), .ZN(n2363) );
  oai22d1 U3854 ( .A1(n2363), .A2(n2362), .B1(n5273), .B2(n2369), .ZN(n4166)
         );
  inv0d0 U3855 ( .I(csrbank6_ien1_w[27]), .ZN(n2364) );
  oai22d1 U3856 ( .A1(n2364), .A2(n2370), .B1(n5275), .B2(n2367), .ZN(n4165)
         );
  inv0d0 U3857 ( .I(csrbank6_ien1_w[28]), .ZN(n2365) );
  oai22d1 U3858 ( .A1(n2365), .A2(n2370), .B1(n5276), .B2(n2367), .ZN(n4164)
         );
  inv0d0 U3859 ( .I(csrbank6_ien1_w[29]), .ZN(n2366) );
  oai22d1 U3860 ( .A1(n2366), .A2(n2370), .B1(n5280), .B2(n2367), .ZN(n4163)
         );
  inv0d0 U3861 ( .I(csrbank6_ien1_w[30]), .ZN(n2368) );
  oai22d1 U3862 ( .A1(n2368), .A2(n2370), .B1(n5283), .B2(n2367), .ZN(n4162)
         );
  inv0d0 U3863 ( .I(csrbank6_ien1_w[31]), .ZN(n2371) );
  oai22d1 U3864 ( .A1(n2371), .A2(n2370), .B1(n5287), .B2(n2369), .ZN(n4161)
         );
  inv0d0 U3865 ( .I(csrbank6_ien2_w[0]), .ZN(n2374) );
  oai21d1 U3866 ( .B1(n2372), .B2(n4959), .A(n5955), .ZN(n2400) );
  nd03d1 U3867 ( .A1(n2373), .A2(n5240), .A3(n5288), .ZN(n2407) );
  buffd1 U3868 ( .I(n2407), .Z(n2404) );
  oai22d1 U3869 ( .A1(n2374), .A2(n2400), .B1(n2472), .B2(n2404), .ZN(n4160)
         );
  inv0d0 U3870 ( .I(csrbank6_ien2_w[1]), .ZN(n2375) );
  oai22d1 U3871 ( .A1(n2375), .A2(n2400), .B1(n2639), .B2(n2404), .ZN(n4159)
         );
  inv0d0 U3872 ( .I(csrbank6_ien2_w[2]), .ZN(n2376) );
  oai22d1 U3873 ( .A1(n2376), .A2(n2400), .B1(n5004), .B2(n2404), .ZN(n4158)
         );
  inv0d0 U3874 ( .I(csrbank6_ien2_w[3]), .ZN(n2377) );
  buffd1 U3875 ( .I(n2625), .Z(n5006) );
  oai22d1 U3876 ( .A1(n2377), .A2(n2400), .B1(n5006), .B2(n2404), .ZN(n4157)
         );
  inv0d0 U3877 ( .I(csrbank6_ien2_w[4]), .ZN(n2378) );
  buffd1 U3878 ( .I(n2400), .Z(n2408) );
  oai22d1 U3879 ( .A1(n2378), .A2(n2408), .B1(n4866), .B2(n2404), .ZN(n4156)
         );
  inv0d0 U3880 ( .I(csrbank6_ien2_w[5]), .ZN(n2379) );
  oai22d1 U3881 ( .A1(n2379), .A2(n2408), .B1(n5010), .B2(n2404), .ZN(n4155)
         );
  inv0d0 U3882 ( .I(csrbank6_ien2_w[6]), .ZN(n2380) );
  oai22d1 U3883 ( .A1(n2380), .A2(n2400), .B1(n5012), .B2(n2404), .ZN(n4154)
         );
  inv0d0 U3884 ( .I(csrbank6_ien2_w[7]), .ZN(n2381) );
  oai22d1 U3885 ( .A1(n2381), .A2(n2400), .B1(n5251), .B2(n2404), .ZN(n4153)
         );
  inv0d0 U3886 ( .I(csrbank6_ien2_w[8]), .ZN(n2382) );
  oai22d1 U3887 ( .A1(n2382), .A2(n2400), .B1(n4783), .B2(n2404), .ZN(n4152)
         );
  inv0d0 U3888 ( .I(csrbank6_ien2_w[9]), .ZN(n2383) );
  oai22d1 U3889 ( .A1(n2383), .A2(n2408), .B1(n5017), .B2(n2404), .ZN(n4151)
         );
  inv0d0 U3890 ( .I(csrbank6_ien2_w[10]), .ZN(n2384) );
  oai22d1 U3891 ( .A1(n2384), .A2(n2400), .B1(n5019), .B2(n2407), .ZN(n4150)
         );
  inv0d0 U3892 ( .I(csrbank6_ien2_w[11]), .ZN(n2385) );
  oai22d1 U3893 ( .A1(n2385), .A2(n2400), .B1(n5254), .B2(n2407), .ZN(n4149)
         );
  inv0d0 U3894 ( .I(csrbank6_ien2_w[12]), .ZN(n2386) );
  oai22d1 U3895 ( .A1(n2386), .A2(n2408), .B1(n5022), .B2(n2407), .ZN(n4148)
         );
  inv0d0 U3896 ( .I(csrbank6_ien2_w[13]), .ZN(n2387) );
  oai22d1 U3897 ( .A1(n2387), .A2(n2400), .B1(n4790), .B2(n2404), .ZN(n4147)
         );
  inv0d0 U3898 ( .I(csrbank6_ien2_w[14]), .ZN(n2388) );
  oai22d1 U3899 ( .A1(n2388), .A2(n2400), .B1(n5026), .B2(n2404), .ZN(n4146)
         );
  inv0d0 U3900 ( .I(csrbank6_ien2_w[15]), .ZN(n2389) );
  oai22d1 U3901 ( .A1(n2389), .A2(n2408), .B1(n4793), .B2(n2407), .ZN(n4145)
         );
  inv0d0 U3902 ( .I(csrbank6_ien2_w[16]), .ZN(n2390) );
  oai22d1 U3903 ( .A1(n2390), .A2(n2408), .B1(n2003), .B2(n2407), .ZN(n4144)
         );
  inv0d0 U3904 ( .I(csrbank6_ien2_w[17]), .ZN(n2391) );
  oai22d1 U3905 ( .A1(n2391), .A2(n2408), .B1(n5259), .B2(n2404), .ZN(n4143)
         );
  inv0d0 U3906 ( .I(csrbank6_ien2_w[18]), .ZN(n2392) );
  oai22d1 U3907 ( .A1(n2392), .A2(n2400), .B1(n5260), .B2(n2404), .ZN(n4142)
         );
  inv0d0 U3908 ( .I(csrbank6_ien2_w[19]), .ZN(n2393) );
  oai22d1 U3909 ( .A1(n2393), .A2(n2408), .B1(n5262), .B2(n2407), .ZN(n4141)
         );
  inv0d0 U3910 ( .I(csrbank6_ien2_w[20]), .ZN(n2394) );
  oai22d1 U3911 ( .A1(n2394), .A2(n2400), .B1(n5263), .B2(n2404), .ZN(n4140)
         );
  inv0d0 U3912 ( .I(csrbank6_ien2_w[21]), .ZN(n2395) );
  oai22d1 U3913 ( .A1(n2395), .A2(n2408), .B1(n5264), .B2(n2407), .ZN(n4139)
         );
  inv0d0 U3914 ( .I(csrbank6_ien2_w[22]), .ZN(n2396) );
  oai22d1 U3915 ( .A1(n2396), .A2(n2400), .B1(n5266), .B2(n2407), .ZN(n4138)
         );
  inv0d0 U3916 ( .I(csrbank6_ien2_w[23]), .ZN(n2397) );
  oai22d1 U3917 ( .A1(n2397), .A2(n2408), .B1(n5268), .B2(n2407), .ZN(n4137)
         );
  inv0d0 U3918 ( .I(csrbank6_ien2_w[24]), .ZN(n2398) );
  oai22d1 U3919 ( .A1(n2398), .A2(n2408), .B1(n5270), .B2(n2407), .ZN(n4136)
         );
  inv0d0 U3920 ( .I(csrbank6_ien2_w[25]), .ZN(n2399) );
  oai22d1 U3921 ( .A1(n2399), .A2(n2408), .B1(n5271), .B2(n2407), .ZN(n4135)
         );
  inv0d0 U3922 ( .I(csrbank6_ien2_w[26]), .ZN(n2401) );
  oai22d1 U3923 ( .A1(n2401), .A2(n2400), .B1(n5273), .B2(n2407), .ZN(n4134)
         );
  inv0d0 U3924 ( .I(csrbank6_ien2_w[27]), .ZN(n2402) );
  oai22d1 U3925 ( .A1(n2402), .A2(n2408), .B1(n5275), .B2(n2407), .ZN(n4133)
         );
  inv0d0 U3926 ( .I(csrbank6_ien2_w[28]), .ZN(n2403) );
  oai22d1 U3927 ( .A1(n2403), .A2(n2408), .B1(n5276), .B2(n2404), .ZN(n4132)
         );
  inv0d0 U3928 ( .I(csrbank6_ien2_w[29]), .ZN(n2405) );
  oai22d1 U3929 ( .A1(n2405), .A2(n2408), .B1(n5280), .B2(n2404), .ZN(n4131)
         );
  inv0d0 U3930 ( .I(csrbank6_ien2_w[30]), .ZN(n2406) );
  oai22d1 U3931 ( .A1(n2406), .A2(n2408), .B1(n5283), .B2(n2407), .ZN(n4130)
         );
  inv0d0 U3932 ( .I(csrbank6_ien2_w[31]), .ZN(n2409) );
  oai22d1 U3933 ( .A1(n2409), .A2(n2408), .B1(n5287), .B2(n2407), .ZN(n4129)
         );
  inv0d0 U3934 ( .I(csrbank6_ien3_w[0]), .ZN(n2411) );
  oaim21d1 U3935 ( .B1(n4683), .B2(n2410), .A(n5340), .ZN(n2435) );
  nd02d1 U3936 ( .A1(n2410), .A2(n4580), .ZN(n2444) );
  buffd1 U3937 ( .I(n2444), .Z(n2437) );
  oai22d1 U3938 ( .A1(n2411), .A2(n2435), .B1(n2472), .B2(n2437), .ZN(n4128)
         );
  inv0d0 U3939 ( .I(csrbank6_ien3_w[1]), .ZN(n2412) );
  oai22d1 U3940 ( .A1(n2412), .A2(n2435), .B1(n4862), .B2(n2437), .ZN(n4127)
         );
  inv0d0 U3941 ( .I(csrbank6_ien3_w[2]), .ZN(n2413) );
  oai22d1 U3942 ( .A1(n2413), .A2(n2435), .B1(n5004), .B2(n2437), .ZN(n4126)
         );
  inv0d0 U3943 ( .I(csrbank6_ien3_w[3]), .ZN(n2414) );
  oai22d1 U3944 ( .A1(n2414), .A2(n2435), .B1(n5006), .B2(n2437), .ZN(n4125)
         );
  inv0d0 U3945 ( .I(csrbank6_ien3_w[4]), .ZN(n2415) );
  buffd1 U3946 ( .I(n2435), .Z(n2445) );
  oai22d1 U3947 ( .A1(n2415), .A2(n2445), .B1(n5008), .B2(n2437), .ZN(n4124)
         );
  inv0d0 U3948 ( .I(csrbank6_ien3_w[5]), .ZN(n2416) );
  oai22d1 U3949 ( .A1(n2416), .A2(n2445), .B1(n5010), .B2(n2437), .ZN(n4123)
         );
  inv0d0 U3950 ( .I(csrbank6_ien3_w[6]), .ZN(n2417) );
  oai22d1 U3951 ( .A1(n2417), .A2(n2445), .B1(n5012), .B2(n2437), .ZN(n4122)
         );
  inv0d0 U3952 ( .I(csrbank6_ien3_w[7]), .ZN(n2418) );
  oai22d1 U3953 ( .A1(n2418), .A2(n2445), .B1(n5251), .B2(n2437), .ZN(n4121)
         );
  inv0d0 U3954 ( .I(csrbank6_ien3_w[8]), .ZN(n2419) );
  oai22d1 U3955 ( .A1(n2419), .A2(n2445), .B1(n5015), .B2(n2437), .ZN(n4120)
         );
  inv0d0 U3956 ( .I(csrbank6_ien3_w[9]), .ZN(n2420) );
  oai22d1 U3957 ( .A1(n2420), .A2(n2435), .B1(n5017), .B2(n2444), .ZN(n4119)
         );
  inv0d0 U3958 ( .I(csrbank6_ien3_w[10]), .ZN(n2421) );
  oai22d1 U3959 ( .A1(n2421), .A2(n2445), .B1(n5019), .B2(n2437), .ZN(n4118)
         );
  inv0d0 U3960 ( .I(csrbank6_ien3_w[11]), .ZN(n2422) );
  oai22d1 U3961 ( .A1(n2422), .A2(n2435), .B1(n4787), .B2(n2437), .ZN(n4117)
         );
  inv0d0 U3962 ( .I(csrbank6_ien3_w[12]), .ZN(n2423) );
  oai22d1 U3963 ( .A1(n2423), .A2(n2445), .B1(n5022), .B2(n2444), .ZN(n4116)
         );
  inv0d0 U3964 ( .I(csrbank6_ien3_w[13]), .ZN(n2424) );
  oai22d1 U3965 ( .A1(n2424), .A2(n2435), .B1(n5024), .B2(n2444), .ZN(n4115)
         );
  inv0d0 U3966 ( .I(csrbank6_ien3_w[14]), .ZN(n2425) );
  oai22d1 U3967 ( .A1(n2425), .A2(n2445), .B1(n5026), .B2(n2444), .ZN(n4114)
         );
  inv0d0 U3968 ( .I(csrbank6_ien3_w[15]), .ZN(n2426) );
  oai22d1 U3969 ( .A1(n2426), .A2(n2435), .B1(n5028), .B2(n2437), .ZN(n4113)
         );
  inv0d0 U3970 ( .I(csrbank6_ien3_w[16]), .ZN(n2427) );
  oai22d1 U3971 ( .A1(n2427), .A2(n2435), .B1(n2003), .B2(n2444), .ZN(n4112)
         );
  inv0d0 U3972 ( .I(csrbank6_ien3_w[17]), .ZN(n2428) );
  oai22d1 U3973 ( .A1(n2428), .A2(n2435), .B1(n5259), .B2(n2437), .ZN(n4111)
         );
  inv0d0 U3974 ( .I(csrbank6_ien3_w[18]), .ZN(n2429) );
  oai22d1 U3975 ( .A1(n2429), .A2(n2445), .B1(n5260), .B2(n2437), .ZN(n4110)
         );
  inv0d0 U3976 ( .I(csrbank6_ien3_w[19]), .ZN(n2430) );
  oai22d1 U3977 ( .A1(n2430), .A2(n2435), .B1(n5262), .B2(n2444), .ZN(n4109)
         );
  inv0d0 U3978 ( .I(csrbank6_ien3_w[20]), .ZN(n2431) );
  oai22d1 U3979 ( .A1(n2431), .A2(n2435), .B1(n5263), .B2(n2444), .ZN(n4108)
         );
  inv0d0 U3980 ( .I(csrbank6_ien3_w[21]), .ZN(n2432) );
  oai22d1 U3981 ( .A1(n2432), .A2(n2435), .B1(n5264), .B2(n2444), .ZN(n4107)
         );
  inv0d0 U3982 ( .I(csrbank6_ien3_w[22]), .ZN(n2433) );
  oai22d1 U3983 ( .A1(n2433), .A2(n2435), .B1(n5266), .B2(n2444), .ZN(n4106)
         );
  inv0d0 U3984 ( .I(csrbank6_ien3_w[23]), .ZN(n2434) );
  oai22d1 U3985 ( .A1(n2434), .A2(n2445), .B1(n5268), .B2(n2437), .ZN(n4105)
         );
  inv0d0 U3986 ( .I(csrbank6_ien3_w[24]), .ZN(n2436) );
  oai22d1 U3987 ( .A1(n2436), .A2(n2435), .B1(n5270), .B2(n2437), .ZN(n4104)
         );
  inv0d0 U3988 ( .I(csrbank6_ien3_w[25]), .ZN(n2438) );
  oai22d1 U3989 ( .A1(n2438), .A2(n2445), .B1(n5271), .B2(n2437), .ZN(n4103)
         );
  inv0d0 U3990 ( .I(csrbank6_ien3_w[26]), .ZN(n2439) );
  oai22d1 U3991 ( .A1(n2439), .A2(n2445), .B1(n5273), .B2(n2444), .ZN(n4102)
         );
  inv0d0 U3992 ( .I(csrbank6_ien3_w[27]), .ZN(n2440) );
  oai22d1 U3993 ( .A1(n2440), .A2(n2445), .B1(n5275), .B2(n2444), .ZN(n4101)
         );
  inv0d0 U3994 ( .I(csrbank6_ien3_w[28]), .ZN(n2441) );
  oai22d1 U3995 ( .A1(n2441), .A2(n2445), .B1(n5276), .B2(n2444), .ZN(n4100)
         );
  inv0d0 U3996 ( .I(csrbank6_ien3_w[29]), .ZN(n2442) );
  oai22d1 U3997 ( .A1(n2442), .A2(n2445), .B1(n5280), .B2(n2444), .ZN(n4099)
         );
  inv0d0 U3998 ( .I(csrbank6_ien3_w[30]), .ZN(n2443) );
  oai22d1 U3999 ( .A1(n2443), .A2(n2445), .B1(n5283), .B2(n2444), .ZN(n4098)
         );
  inv0d0 U4000 ( .I(csrbank6_ien3_w[31]), .ZN(n2446) );
  oai22d1 U4001 ( .A1(n2446), .A2(n2445), .B1(n5287), .B2(n2444), .ZN(n4097)
         );
  nd02d0 U4002 ( .A1(n2647), .A2(n2450), .ZN(n2448) );
  oai21d1 U4003 ( .B1(n2448), .B2(n5000), .A(n2447), .ZN(n4096) );
  nd02d0 U4004 ( .A1(n2450), .A2(n2449), .ZN(n2461) );
  oai21d1 U4005 ( .B1(csrbank5_oe0_w), .B2(n2453), .A(n5955), .ZN(n2452) );
  aoi21d1 U4006 ( .B1(n2453), .B2(n4808), .A(n2452), .ZN(n4095) );
  nr02d0 U4007 ( .A1(n2454), .A2(n2461), .ZN(n2456) );
  oai21d1 U4008 ( .B1(csrbank5_ien0_w), .B2(n2456), .A(n5955), .ZN(n2455) );
  aoi21d1 U4009 ( .B1(n2456), .B2(n5290), .A(n2455), .ZN(n4094) );
  inv0d0 U4010 ( .I(n2457), .ZN(n2458) );
  nr02d0 U4011 ( .A1(n2458), .A2(n2461), .ZN(n2460) );
  oai21d1 U4012 ( .B1(gpio_mode0_pad), .B2(n2460), .A(n5319), .ZN(n2459) );
  aoi21d1 U4013 ( .B1(n2460), .B2(n266), .A(n2459), .ZN(n4093) );
  nr02d0 U4014 ( .A1(n2462), .A2(n2461), .ZN(n2464) );
  oai21d1 U4015 ( .B1(gpio_mode1_pad), .B2(n2464), .A(n5955), .ZN(n2463) );
  aoi21d1 U4016 ( .B1(n2464), .B2(n2472), .A(n2463), .ZN(n4092) );
  nd03d0 U4017 ( .A1(n2468), .A2(uart_enabled_o), .A3(n5956), .ZN(n2467) );
  oai21d1 U4018 ( .B1(n2468), .B2(n4955), .A(n2467), .ZN(n4091) );
  nr04d0 U4019 ( .A1(n4811), .A2(n3060), .A3(n2470), .A4(n2469), .ZN(n2473) );
  oai21d1 U4020 ( .B1(debug_mode), .B2(n2473), .A(n5319), .ZN(n2471) );
  aoi21d1 U4021 ( .B1(n2473), .B2(n5290), .A(n2471), .ZN(n4090) );
  nd03d0 U4022 ( .A1(n2478), .A2(debug_oeb), .A3(n5340), .ZN(n2477) );
  oai21d1 U4023 ( .B1(n2478), .B2(n4955), .A(n2477), .ZN(n4089) );
  nr02d0 U4024 ( .A1(n2479), .A2(dbg_uart_count[15]), .ZN(n2489) );
  nd12d0 U4025 ( .A1(dbg_uart_count[16]), .A2(n2489), .ZN(n2487) );
  nr02d0 U4026 ( .A1(n2487), .A2(dbg_uart_count[17]), .ZN(n2484) );
  inv0d0 U4027 ( .I(n2484), .ZN(n2480) );
  oai21d1 U4028 ( .B1(dbg_uart_count[18]), .B2(n2480), .A(dbg_uart_count[19]), 
        .ZN(n2481) );
  inv0d0 U4029 ( .I(n2481), .ZN(n2483) );
  nr02d0 U4030 ( .A1(n2482), .A2(n5492), .ZN(n5318) );
  nd12d0 U4031 ( .A1(n2483), .A2(n5318), .ZN(n4087) );
  aoim22d1 U4032 ( .A1(dbg_uart_count[18]), .A2(n2484), .B1(n2484), .B2(
        dbg_uart_count[18]), .Z(n2485) );
  oaim21d1 U4033 ( .B1(n2485), .B2(n2497), .A(n5318), .ZN(n4086) );
  inv0d0 U4034 ( .I(dbg_uart_count[17]), .ZN(n2486) );
  aoim22d1 U4035 ( .A1(n2487), .A2(n2486), .B1(n2486), .B2(n2487), .Z(n2488)
         );
  oaim21d1 U4036 ( .B1(n2488), .B2(n2497), .A(n5318), .ZN(n4085) );
  aoim22d1 U4037 ( .A1(dbg_uart_count[16]), .A2(n2489), .B1(n2489), .B2(
        dbg_uart_count[16]), .Z(n2490) );
  oaim21d1 U4038 ( .B1(n2490), .B2(n2497), .A(n5318), .ZN(n4084) );
  aoim22d1 U4039 ( .A1(dbg_uart_count[14]), .A2(n2491), .B1(n2491), .B2(
        dbg_uart_count[14]), .Z(n2492) );
  oaim21d1 U4040 ( .B1(n2492), .B2(n2497), .A(n5318), .ZN(n4082) );
  inv0d0 U4041 ( .I(n2493), .ZN(n2494) );
  aoim22d1 U4042 ( .A1(dbg_uart_count[9]), .A2(n2494), .B1(n2494), .B2(
        dbg_uart_count[9]), .Z(n2495) );
  oaim21d1 U4043 ( .B1(n2495), .B2(n2497), .A(n5318), .ZN(n4077) );
  aoim22d1 U4044 ( .A1(dbg_uart_count[6]), .A2(n2496), .B1(n2496), .B2(
        dbg_uart_count[6]), .Z(n2498) );
  oaim21d1 U4045 ( .B1(n2498), .B2(n2497), .A(n5318), .ZN(n4074) );
  aoi21d1 U4046 ( .B1(dbg_uart_cmd[0]), .B2(dbg_uart_cmd[1]), .A(
        dbg_uart_cmd[2]), .ZN(n2499) );
  oai211d1 U4047 ( .C1(dbg_uart_cmd[0]), .C2(dbg_uart_cmd[1]), .A(n2501), .B(
        n2499), .ZN(n2507) );
  inv0d0 U4048 ( .I(n2500), .ZN(n2503) );
  nd03d0 U4049 ( .A1(n2501), .A2(dbg_uart_cmd[1]), .A3(n5960), .ZN(n2502) );
  aon211d1 U4050 ( .C1(n2503), .C2(n2502), .B(n2506), .A(dbg_uart_incr), .ZN(
        n2505) );
  oan211d1 U4051 ( .C1(n2507), .C2(n2506), .B(n2505), .A(n2504), .ZN(n4068) );
  inv0d0 U4052 ( .I(n5300), .ZN(n5989) );
  nd02d1 U4053 ( .A1(n5989), .A2(n2508), .ZN(n6019) );
  aon211d1 U4054 ( .C1(dbg_uart_tx_tick), .C2(dbg_uart_tx_data[0]), .B(n5990), 
        .A(n6019), .ZN(n2509) );
  oai31d1 U4055 ( .B1(dbg_uart_tx_tick), .B2(n5990), .B3(n2510), .A(n2509), 
        .ZN(n4067) );
  inv0d0 U4056 ( .I(uart_rx_fifo_rdport_adr[0]), .ZN(n3042) );
  inv0d0 U4057 ( .I(n3022), .ZN(n2517) );
  aoi211d1 U4058 ( .C1(n3020), .C2(n3042), .A(n5111), .B(n2517), .ZN(n4066) );
  nr02d0 U4059 ( .A1(n2511), .A2(n3022), .ZN(n2513) );
  aoi211d1 U4060 ( .C1(n2511), .C2(n3022), .A(n4878), .B(n2513), .ZN(n4065) );
  nr02d0 U4061 ( .A1(n2512), .A2(n3022), .ZN(n2514) );
  aoim211d1 U4062 ( .C1(uart_rx_fifo_rdport_adr[2]), .C2(n2513), .A(n5111), 
        .B(n2514), .ZN(n4064) );
  nr02d0 U4063 ( .A1(uart_rx_fifo_rdport_adr[3]), .A2(n2514), .ZN(n2515) );
  aoi211d1 U4064 ( .C1(n3033), .C2(n2517), .A(n2516), .B(n2515), .ZN(n4063) );
  nd03d0 U4065 ( .A1(uart_phy_rx_rx), .A2(n2519), .A3(n2518), .ZN(n2532) );
  inv0d0 U4066 ( .I(uart_rx_fifo_produce[0]), .ZN(n2913) );
  nr02d0 U4067 ( .A1(n2532), .A2(n2913), .ZN(n2909) );
  aoi211d1 U4068 ( .C1(n2532), .C2(n2913), .A(n5492), .B(n2909), .ZN(n4062) );
  inv0d0 U4069 ( .I(uart_rx_fifo_produce[1]), .ZN(n2901) );
  inv0d0 U4070 ( .I(n2909), .ZN(n2520) );
  aoi221d1 U4071 ( .B1(uart_rx_fifo_produce[1]), .B2(n2909), .C1(n2901), .C2(
        n2520), .A(n5492), .ZN(n4061) );
  inv0d0 U4072 ( .I(uart_rx_fifo_produce[2]), .ZN(n2902) );
  nd02d0 U4073 ( .A1(uart_rx_fifo_produce[1]), .A2(n2909), .ZN(n2521) );
  nd02d0 U4074 ( .A1(uart_rx_fifo_produce[2]), .A2(uart_rx_fifo_produce[1]), 
        .ZN(n2916) );
  nr02d0 U4075 ( .A1(n2916), .A2(n2520), .ZN(n2522) );
  aoi211d1 U4076 ( .C1(n2902), .C2(n2521), .A(n2516), .B(n2522), .ZN(n4060) );
  nd02d0 U4077 ( .A1(uart_rx_fifo_produce[3]), .A2(n2909), .ZN(n2903) );
  nr02d1 U4078 ( .A1(n2916), .A2(n2903), .ZN(n2893) );
  aoim211d1 U4079 ( .C1(uart_rx_fifo_produce[3]), .C2(n2522), .A(n5100), .B(
        n2893), .ZN(n4059) );
  inv0d0 U4080 ( .I(n2532), .ZN(n2915) );
  nr02d0 U4081 ( .A1(n2915), .A2(n3020), .ZN(n2543) );
  nr02d0 U4082 ( .A1(n3046), .A2(n2532), .ZN(n2544) );
  nr02d0 U4083 ( .A1(n2543), .A2(n2544), .ZN(n2547) );
  nd02d0 U4084 ( .A1(n2547), .A2(n5301), .ZN(n2537) );
  or02d0 U4085 ( .A1(n2547), .A2(n5111), .Z(n2539) );
  inv0d0 U4086 ( .I(uart_rx_fifo_level0[0]), .ZN(n2523) );
  aoi22d1 U4087 ( .A1(uart_rx_fifo_level0[0]), .A2(n2537), .B1(n2539), .B2(
        n2523), .ZN(n4058) );
  inv0d0 U4088 ( .I(uart_rx_fifo_level0[3]), .ZN(n2524) );
  nd04d0 U4089 ( .A1(uart_rx_fifo_level0[2]), .A2(uart_rx_fifo_level0[1]), 
        .A3(uart_rx_fifo_level0[0]), .A4(n2915), .ZN(n2535) );
  nr02d0 U4090 ( .A1(n2524), .A2(n2535), .ZN(n2526) );
  oan211d1 U4091 ( .C1(n2526), .C2(n2550), .B(uart_rx_fifo_level0[4]), .A(
        n2539), .ZN(n2525) );
  oai21d1 U4092 ( .B1(n2526), .B2(uart_rx_fifo_level0[4]), .A(n2525), .ZN(
        n2527) );
  oai21d1 U4093 ( .B1(n2537), .B2(n2549), .A(n2527), .ZN(n4057) );
  nr03d0 U4094 ( .A1(uart_rx_fifo_level0[2]), .A2(uart_rx_fifo_level0[1]), 
        .A3(uart_rx_fifo_level0[0]), .ZN(n2528) );
  nd02d0 U4095 ( .A1(n2528), .A2(n2543), .ZN(n2533) );
  aoi21d1 U4096 ( .B1(n2535), .B2(n2533), .A(n2547), .ZN(n2530) );
  oai21d1 U4097 ( .B1(uart_rx_fifo_level0[3]), .B2(n2530), .A(n5319), .ZN(
        n2529) );
  aoi21d1 U4098 ( .B1(uart_rx_fifo_level0[3]), .B2(n2530), .A(n2529), .ZN(
        n4056) );
  nr02d0 U4099 ( .A1(uart_rx_fifo_level0[1]), .A2(uart_rx_fifo_level0[0]), 
        .ZN(n2541) );
  inv0d0 U4100 ( .I(uart_rx_fifo_level0[2]), .ZN(n2538) );
  nd03d0 U4101 ( .A1(uart_rx_fifo_level0[1]), .A2(uart_rx_fifo_level0[0]), 
        .A3(n2915), .ZN(n2531) );
  aoi22d1 U4102 ( .A1(n2541), .A2(n2532), .B1(n2538), .B2(n2531), .ZN(n2536)
         );
  inv0d0 U4103 ( .I(n2533), .ZN(n2534) );
  aoi21d1 U4104 ( .B1(n2536), .B2(n2535), .A(n2534), .ZN(n2540) );
  oai22d1 U4105 ( .A1(n2540), .A2(n2539), .B1(n2538), .B2(n2537), .ZN(n4055)
         );
  inv0d0 U4106 ( .I(uart_rx_fifo_level0[1]), .ZN(n2546) );
  aoi21d1 U4107 ( .B1(uart_rx_fifo_level0[0]), .B2(uart_rx_fifo_level0[1]), 
        .A(n2541), .ZN(n2542) );
  mx02d1 U4108 ( .I0(n2544), .I1(n2543), .S(n2542), .Z(n2545) );
  aoi211d1 U4109 ( .C1(n2547), .C2(n2546), .A(n4878), .B(n2545), .ZN(n4054) );
  aoi31d1 U4110 ( .B1(n2550), .B2(n2549), .B3(n2548), .A(sys_rst), .ZN(n4053)
         );
  nd02d0 U4111 ( .A1(uart_phy_tx_tick), .A2(uart_phy_tx_count[0]), .ZN(n2669)
         );
  inv0d0 U4112 ( .I(uart_phy_tx_count[2]), .ZN(n2671) );
  nd02d0 U4113 ( .A1(rs232phy_rs232phytx_state), .A2(n2671), .ZN(n2552) );
  inv0d0 U4114 ( .I(uart_phy_tx_count[3]), .ZN(n2551) );
  nr04d0 U4115 ( .A1(uart_phy_tx_count[1]), .A2(n2669), .A3(n2552), .A4(n2551), 
        .ZN(n2665) );
  nr02d0 U4116 ( .A1(n2665), .A2(n2666), .ZN(n2644) );
  inv0d0 U4117 ( .I(uart_tx_fifo_level0[4]), .ZN(n2567) );
  an02d0 U4118 ( .A1(n2567), .A2(n2563), .Z(n2646) );
  nr02d1 U4119 ( .A1(n2644), .A2(n2646), .ZN(n2845) );
  inv0d0 U4120 ( .I(n2845), .ZN(n2809) );
  inv0d0 U4121 ( .I(uart_tx_fifo_rdport_adr[0]), .ZN(n2806) );
  nr02d0 U4122 ( .A1(n2809), .A2(n2806), .ZN(n2767) );
  aoi211d1 U4123 ( .C1(n2809), .C2(n2806), .A(n4878), .B(n2767), .ZN(n4052) );
  nd02d0 U4124 ( .A1(uart_tx_fifo_rdport_adr[1]), .A2(n2767), .ZN(n2553) );
  ora211d1 U4125 ( .C1(uart_tx_fifo_rdport_adr[1]), .C2(n2767), .A(n5956), .B(
        n2553), .Z(n4051) );
  inv0d0 U4126 ( .I(uart_tx_fifo_rdport_adr[2]), .ZN(n2677) );
  nr02d0 U4127 ( .A1(n2677), .A2(n2553), .ZN(n2554) );
  aoi211d1 U4128 ( .C1(n2677), .C2(n2553), .A(sys_rst), .B(n2554), .ZN(n4050)
         );
  inv0d0 U4129 ( .I(uart_tx_fifo_rdport_adr[1]), .ZN(n2674) );
  inv0d0 U4130 ( .I(uart_tx_fifo_rdport_adr[3]), .ZN(n2680) );
  nr03d1 U4131 ( .A1(n2677), .A2(n2674), .A3(n2680), .ZN(n2801) );
  nr02d0 U4132 ( .A1(n2554), .A2(uart_tx_fifo_rdport_adr[3]), .ZN(n2555) );
  aoi211d1 U4133 ( .C1(n2767), .C2(n2801), .A(n5111), .B(n2555), .ZN(n4049) );
  nd03d1 U4134 ( .A1(n4683), .A2(n2557), .A3(n2556), .ZN(n2594) );
  inv0d0 U4135 ( .I(uart_tx_fifo_produce[0]), .ZN(n2613) );
  aoi211d1 U4136 ( .C1(n2594), .C2(n2613), .A(sys_rst), .B(n2621), .ZN(n4048)
         );
  inv0d0 U4137 ( .I(uart_tx_fifo_produce[1]), .ZN(n2615) );
  inv0d0 U4138 ( .I(n2621), .ZN(n2558) );
  aoi211d1 U4139 ( .C1(n2615), .C2(n2558), .A(n4878), .B(n2559), .ZN(n4047) );
  inv0d0 U4140 ( .I(n2591), .ZN(n2560) );
  aoim211d1 U4141 ( .C1(uart_tx_fifo_produce[2]), .C2(n2559), .A(n5111), .B(
        n2560), .ZN(n4046) );
  inv0d0 U4142 ( .I(uart_tx_fifo_produce[3]), .ZN(n2620) );
  oan211d1 U4143 ( .C1(n2560), .C2(n2620), .B(n2611), .A(n5492), .ZN(n4045) );
  nd02d0 U4144 ( .A1(n2845), .A2(n2594), .ZN(n2574) );
  oai21d1 U4145 ( .B1(n2845), .B2(n2594), .A(n2574), .ZN(n2589) );
  inv0d0 U4146 ( .I(n2589), .ZN(n2562) );
  aoi221d1 U4147 ( .B1(uart_tx_fifo_level0[0]), .B2(n2589), .C1(n2561), .C2(
        n2562), .A(sys_rst), .ZN(n4044) );
  nd02d0 U4148 ( .A1(n2562), .A2(n5956), .ZN(n2579) );
  inv0d0 U4149 ( .I(uart_tx_fifo_level0[3]), .ZN(n2570) );
  nd02d0 U4150 ( .A1(uart_tx_fifo_level0[1]), .A2(uart_tx_fifo_level0[0]), 
        .ZN(n2575) );
  nr04d0 U4151 ( .A1(n2580), .A2(n2570), .A3(n2594), .A4(n2575), .ZN(n2565) );
  nd02d0 U4152 ( .A1(n5955), .A2(n2589), .ZN(n2581) );
  oan211d1 U4153 ( .C1(n2565), .C2(n2563), .B(uart_tx_fifo_level0[4]), .A(
        n2581), .ZN(n2564) );
  oai21d1 U4154 ( .B1(n2565), .B2(uart_tx_fifo_level0[4]), .A(n2564), .ZN(
        n2566) );
  oai21d1 U4155 ( .B1(n2579), .B2(n2567), .A(n2566), .ZN(n4043) );
  nr02d0 U4156 ( .A1(n2569), .A2(n2574), .ZN(n2577) );
  nr03d0 U4157 ( .A1(n2580), .A2(n2594), .A3(n2575), .ZN(n2573) );
  inv0d0 U4158 ( .I(n2574), .ZN(n2587) );
  aoi31d1 U4159 ( .B1(uart_tx_fifo_level0[2]), .B2(uart_tx_fifo_level0[1]), 
        .B3(uart_tx_fifo_level0[0]), .A(n2594), .ZN(n2568) );
  aoi211d1 U4160 ( .C1(n2587), .C2(n2569), .A(n2568), .B(n2570), .ZN(n2571) );
  oai22d1 U4161 ( .A1(n2571), .A2(n2581), .B1(n2570), .B2(n2579), .ZN(n2572)
         );
  ora31d1 U4162 ( .B1(uart_tx_fifo_level0[3]), .B2(n2577), .B3(n2573), .A(
        n2572), .Z(n4042) );
  nr02d0 U4163 ( .A1(uart_tx_fifo_level0[1]), .A2(uart_tx_fifo_level0[0]), 
        .ZN(n2584) );
  inv0d0 U4164 ( .I(n2575), .ZN(n2583) );
  oai22d1 U4165 ( .A1(n2584), .A2(n2574), .B1(n2583), .B2(n2594), .ZN(n2578)
         );
  nr03d0 U4166 ( .A1(uart_tx_fifo_level0[2]), .A2(n2594), .A3(n2575), .ZN(
        n2576) );
  aoi211d1 U4167 ( .C1(uart_tx_fifo_level0[2]), .C2(n2578), .A(n2577), .B(
        n2576), .ZN(n2582) );
  oai22d1 U4168 ( .A1(n2582), .A2(n2581), .B1(n2580), .B2(n2579), .ZN(n4041)
         );
  oai21d1 U4169 ( .B1(n2594), .B2(n2845), .A(n2586), .ZN(n2585) );
  oai21d1 U4170 ( .B1(n2587), .B2(n2586), .A(n2585), .ZN(n2588) );
  oan211d1 U4171 ( .C1(n2590), .C2(n2589), .B(n2588), .A(n4878), .ZN(n4040) );
  nr02d1 U4172 ( .A1(n2620), .A2(n2591), .ZN(n2593) );
  inv0d0 U4173 ( .I(\storage[15][0] ), .ZN(n2682) );
  inv0d0 U4174 ( .I(n2593), .ZN(n2592) );
  aoi22d1 U4175 ( .A1(n2593), .A2(n266), .B1(n2682), .B2(n2592), .ZN(n4039) );
  inv0d0 U4176 ( .I(\storage[15][1] ), .ZN(n2814) );
  aoi22d1 U4177 ( .A1(n2593), .A2(n2639), .B1(n2814), .B2(n2592), .ZN(n4038)
         );
  aoim22d1 U4178 ( .A1(n2593), .A2(n5004), .B1(\storage[15][2] ), .B2(n2593), 
        .Z(n4037) );
  aoim22d1 U4179 ( .A1(n2593), .A2(n5246), .B1(\storage[15][3] ), .B2(n2593), 
        .Z(n4036) );
  aoim22d1 U4180 ( .A1(n2593), .A2(n5247), .B1(\storage[15][4] ), .B2(n2593), 
        .Z(n4035) );
  inv0d0 U4181 ( .I(\storage[15][5] ), .ZN(n2749) );
  aoi22d1 U4182 ( .A1(n2593), .A2(n2640), .B1(n2749), .B2(n2592), .ZN(n4034)
         );
  inv0d0 U4183 ( .I(\storage[15][6] ), .ZN(n2723) );
  aoi22d1 U4184 ( .A1(n2593), .A2(n5249), .B1(n2723), .B2(n2592), .ZN(n4033)
         );
  inv0d0 U4185 ( .I(\storage[15][7] ), .ZN(n2695) );
  aoi22d1 U4186 ( .A1(n2593), .A2(n3071), .B1(n2695), .B2(n2592), .ZN(n4032)
         );
  inv0d0 U4187 ( .I(uart_tx_fifo_produce[2]), .ZN(n2616) );
  inv0d0 U4188 ( .I(n2594), .ZN(n2614) );
  aoim22d1 U4189 ( .A1(n2596), .A2(n5290), .B1(\storage[14][0] ), .B2(n2596), 
        .Z(n4031) );
  inv0d0 U4190 ( .I(\storage[14][1] ), .ZN(n2834) );
  inv0d0 U4191 ( .I(n2596), .ZN(n2595) );
  aoi22d1 U4192 ( .A1(n2596), .A2(n4862), .B1(n2834), .B2(n2595), .ZN(n4030)
         );
  aoim22d1 U4193 ( .A1(n2596), .A2(n5004), .B1(\storage[14][2] ), .B2(n2596), 
        .Z(n4029) );
  aoim22d1 U4194 ( .A1(n2596), .A2(n5006), .B1(\storage[14][3] ), .B2(n2596), 
        .Z(n4028) );
  aoim22d1 U4195 ( .A1(n2596), .A2(n5008), .B1(\storage[14][4] ), .B2(n2596), 
        .Z(n4027) );
  aoim22d1 U4196 ( .A1(n2596), .A2(n5010), .B1(\storage[14][5] ), .B2(n2596), 
        .Z(n4026) );
  inv0d0 U4197 ( .I(\storage[14][6] ), .ZN(n2735) );
  aoi22d1 U4198 ( .A1(n2596), .A2(n5012), .B1(n2735), .B2(n2595), .ZN(n4025)
         );
  inv0d0 U4199 ( .I(\storage[14][7] ), .ZN(n2714) );
  aoi22d1 U4200 ( .A1(n2596), .A2(n3071), .B1(n2714), .B2(n2595), .ZN(n4024)
         );
  nr02d1 U4201 ( .A1(n2624), .A2(n2605), .ZN(n2598) );
  aoim22d1 U4202 ( .A1(n2598), .A2(n4808), .B1(\storage[13][0] ), .B2(n2598), 
        .Z(n4023) );
  inv0d0 U4203 ( .I(\storage[13][1] ), .ZN(n2817) );
  inv0d0 U4204 ( .I(n2598), .ZN(n2597) );
  aoi22d1 U4205 ( .A1(n2598), .A2(n4862), .B1(n2817), .B2(n2597), .ZN(n4022)
         );
  aoim22d1 U4206 ( .A1(n2598), .A2(n5004), .B1(\storage[13][2] ), .B2(n2598), 
        .Z(n4021) );
  aoim22d1 U4207 ( .A1(n2598), .A2(n5006), .B1(\storage[13][3] ), .B2(n2598), 
        .Z(n4020) );
  aoim22d1 U4208 ( .A1(n2598), .A2(n5008), .B1(\storage[13][4] ), .B2(n2598), 
        .Z(n4019) );
  inv0d0 U4209 ( .I(\storage[13][5] ), .ZN(n2755) );
  aoi22d1 U4210 ( .A1(n2598), .A2(n5248), .B1(n2755), .B2(n2597), .ZN(n4018)
         );
  inv0d0 U4211 ( .I(\storage[13][6] ), .ZN(n2722) );
  aoi22d1 U4212 ( .A1(n2598), .A2(n2641), .B1(n2722), .B2(n2597), .ZN(n4017)
         );
  inv0d0 U4213 ( .I(\storage[13][7] ), .ZN(n2701) );
  aoi22d1 U4214 ( .A1(n2598), .A2(n3071), .B1(n2701), .B2(n2597), .ZN(n4016)
         );
  nr02d1 U4215 ( .A1(n2608), .A2(n2624), .ZN(n2600) );
  aoim22d1 U4216 ( .A1(n2600), .A2(n266), .B1(\storage[12][0] ), .B2(n2600), 
        .Z(n4015) );
  inv0d0 U4217 ( .I(\storage[12][1] ), .ZN(n2838) );
  inv0d0 U4218 ( .I(n2600), .ZN(n2599) );
  aoi22d1 U4219 ( .A1(n2600), .A2(n4862), .B1(n2838), .B2(n2599), .ZN(n4014)
         );
  aoim22d1 U4220 ( .A1(n2600), .A2(n5004), .B1(\storage[12][2] ), .B2(n2600), 
        .Z(n4013) );
  aoim22d1 U4221 ( .A1(n2600), .A2(n5246), .B1(\storage[12][3] ), .B2(n2600), 
        .Z(n4012) );
  aoim22d1 U4222 ( .A1(n2600), .A2(n5247), .B1(\storage[12][4] ), .B2(n2600), 
        .Z(n4011) );
  aoim22d1 U4223 ( .A1(n2600), .A2(n5248), .B1(\storage[12][5] ), .B2(n2600), 
        .Z(n4010) );
  inv0d0 U4224 ( .I(\storage[12][6] ), .ZN(n2739) );
  aoi22d1 U4225 ( .A1(n2600), .A2(n2641), .B1(n2739), .B2(n2599), .ZN(n4009)
         );
  inv0d0 U4226 ( .I(\storage[12][7] ), .ZN(n2708) );
  aoi22d1 U4227 ( .A1(n2600), .A2(n3071), .B1(n2708), .B2(n2599), .ZN(n4008)
         );
  nd02d0 U4228 ( .A1(uart_tx_fifo_produce[1]), .A2(n2616), .ZN(n2630) );
  nr02d1 U4229 ( .A1(n2605), .A2(n2630), .ZN(n2602) );
  inv0d0 U4230 ( .I(\storage[11][0] ), .ZN(n2676) );
  inv0d0 U4231 ( .I(n2602), .ZN(n2601) );
  aoi22d1 U4232 ( .A1(n2602), .A2(n4808), .B1(n2676), .B2(n2601), .ZN(n4007)
         );
  inv0d0 U4233 ( .I(\storage[11][1] ), .ZN(n2812) );
  aoi22d1 U4234 ( .A1(n2602), .A2(n2639), .B1(n2812), .B2(n2601), .ZN(n4006)
         );
  aoim22d1 U4235 ( .A1(n2602), .A2(n5004), .B1(\storage[11][2] ), .B2(n2602), 
        .Z(n4005) );
  aoim22d1 U4236 ( .A1(n2602), .A2(n5006), .B1(\storage[11][3] ), .B2(n2602), 
        .Z(n4004) );
  aoim22d1 U4237 ( .A1(n2602), .A2(n5008), .B1(\storage[11][4] ), .B2(n2602), 
        .Z(n4003) );
  inv0d0 U4238 ( .I(\storage[11][5] ), .ZN(n2750) );
  aoi22d1 U4239 ( .A1(n2602), .A2(n2640), .B1(n2750), .B2(n2601), .ZN(n4002)
         );
  inv0d0 U4240 ( .I(\storage[11][6] ), .ZN(n2725) );
  aoi22d1 U4241 ( .A1(n2602), .A2(n5249), .B1(n2725), .B2(n2601), .ZN(n4001)
         );
  inv0d0 U4242 ( .I(\storage[11][7] ), .ZN(n2694) );
  aoi22d1 U4243 ( .A1(n2602), .A2(n3071), .B1(n2694), .B2(n2601), .ZN(n4000)
         );
  nr02d1 U4244 ( .A1(n2608), .A2(n2630), .ZN(n2604) );
  aoim22d1 U4245 ( .A1(n2604), .A2(n5290), .B1(\storage[10][0] ), .B2(n2604), 
        .Z(n3999) );
  inv0d0 U4246 ( .I(\storage[10][1] ), .ZN(n2826) );
  inv0d0 U4247 ( .I(n2604), .ZN(n2603) );
  aoi22d1 U4248 ( .A1(n2604), .A2(n4862), .B1(n2826), .B2(n2603), .ZN(n3998)
         );
  aoim22d1 U4249 ( .A1(n2604), .A2(n5004), .B1(\storage[10][2] ), .B2(n2604), 
        .Z(n3997) );
  aoim22d1 U4250 ( .A1(n2604), .A2(n2625), .B1(\storage[10][3] ), .B2(n2604), 
        .Z(n3996) );
  aoim22d1 U4251 ( .A1(n2604), .A2(n4866), .B1(\storage[10][4] ), .B2(n2604), 
        .Z(n3995) );
  aoim22d1 U4252 ( .A1(n2604), .A2(n5010), .B1(\storage[10][5] ), .B2(n2604), 
        .Z(n3994) );
  inv0d0 U4253 ( .I(\storage[10][6] ), .ZN(n2741) );
  aoi22d1 U4254 ( .A1(n2604), .A2(n2641), .B1(n2741), .B2(n2603), .ZN(n3993)
         );
  inv0d0 U4255 ( .I(\storage[10][7] ), .ZN(n2707) );
  aoi22d1 U4256 ( .A1(n2604), .A2(n3071), .B1(n2707), .B2(n2603), .ZN(n3992)
         );
  nd02d0 U4257 ( .A1(n2616), .A2(n2615), .ZN(n2638) );
  nr02d1 U4258 ( .A1(n2605), .A2(n2638), .ZN(n2607) );
  inv0d0 U4259 ( .I(\storage[9][0] ), .ZN(n2681) );
  inv0d0 U4260 ( .I(n2607), .ZN(n2606) );
  aoi22d1 U4261 ( .A1(n2607), .A2(n5290), .B1(n2681), .B2(n2606), .ZN(n3991)
         );
  inv0d0 U4262 ( .I(\storage[9][1] ), .ZN(n2816) );
  aoi22d1 U4263 ( .A1(n2607), .A2(n5294), .B1(n2816), .B2(n2606), .ZN(n3990)
         );
  aoim22d1 U4264 ( .A1(n2607), .A2(n5004), .B1(\storage[9][2] ), .B2(n2607), 
        .Z(n3989) );
  aoim22d1 U4265 ( .A1(n2607), .A2(n2625), .B1(\storage[9][3] ), .B2(n2607), 
        .Z(n3988) );
  aoim22d1 U4266 ( .A1(n2607), .A2(n4866), .B1(\storage[9][4] ), .B2(n2607), 
        .Z(n3987) );
  inv0d0 U4267 ( .I(\storage[9][5] ), .ZN(n2754) );
  aoi22d1 U4268 ( .A1(n2607), .A2(n2640), .B1(n2754), .B2(n2606), .ZN(n3986)
         );
  inv0d0 U4269 ( .I(\storage[9][6] ), .ZN(n2726) );
  aoi22d1 U4270 ( .A1(n2607), .A2(n2641), .B1(n2726), .B2(n2606), .ZN(n3985)
         );
  inv0d0 U4271 ( .I(\storage[9][7] ), .ZN(n2697) );
  aoi22d1 U4272 ( .A1(n2607), .A2(n3071), .B1(n2697), .B2(n2606), .ZN(n3984)
         );
  nr02d1 U4273 ( .A1(n2608), .A2(n2638), .ZN(n2610) );
  aoim22d1 U4274 ( .A1(n2610), .A2(n4808), .B1(\storage[8][0] ), .B2(n2610), 
        .Z(n3983) );
  inv0d0 U4275 ( .I(\storage[8][1] ), .ZN(n2830) );
  inv0d0 U4276 ( .I(n2610), .ZN(n2609) );
  aoi22d1 U4277 ( .A1(n2610), .A2(n4862), .B1(n2830), .B2(n2609), .ZN(n3982)
         );
  aoim22d1 U4278 ( .A1(n2610), .A2(n5004), .B1(\storage[8][2] ), .B2(n2610), 
        .Z(n3981) );
  aoim22d1 U4279 ( .A1(n2610), .A2(n5246), .B1(\storage[8][3] ), .B2(n2610), 
        .Z(n3980) );
  aoim22d1 U4280 ( .A1(n2610), .A2(n5247), .B1(\storage[8][4] ), .B2(n2610), 
        .Z(n3979) );
  aoim22d1 U4281 ( .A1(n2610), .A2(n5248), .B1(\storage[8][5] ), .B2(n2610), 
        .Z(n3978) );
  inv0d0 U4282 ( .I(\storage[8][6] ), .ZN(n2740) );
  aoi22d1 U4283 ( .A1(n2610), .A2(n5012), .B1(n2740), .B2(n2609), .ZN(n3977)
         );
  inv0d0 U4284 ( .I(\storage[8][7] ), .ZN(n2710) );
  aoi22d1 U4285 ( .A1(n2610), .A2(n3071), .B1(n2710), .B2(n2609), .ZN(n3976)
         );
  inv0d1 U4286 ( .I(n2611), .ZN(n2612) );
  aoim22d1 U4287 ( .A1(n2612), .A2(n4808), .B1(\storage[7][0] ), .B2(n2612), 
        .Z(n3975) );
  inv0d0 U4288 ( .I(\storage[7][1] ), .ZN(n2818) );
  aoi22d1 U4289 ( .A1(n2612), .A2(n5294), .B1(n2818), .B2(n2611), .ZN(n3974)
         );
  aoim22d1 U4290 ( .A1(n2612), .A2(n5004), .B1(\storage[7][2] ), .B2(n2612), 
        .Z(n3973) );
  aoim22d1 U4291 ( .A1(n2612), .A2(n5006), .B1(\storage[7][3] ), .B2(n2612), 
        .Z(n3972) );
  aoim22d1 U4292 ( .A1(n2612), .A2(n5008), .B1(\storage[7][4] ), .B2(n2612), 
        .Z(n3971) );
  inv0d0 U4293 ( .I(\storage[7][5] ), .ZN(n2751) );
  aoi22d1 U4294 ( .A1(n2612), .A2(n2640), .B1(n2751), .B2(n2611), .ZN(n3970)
         );
  inv0d0 U4295 ( .I(\storage[7][6] ), .ZN(n2727) );
  aoi22d1 U4296 ( .A1(n2612), .A2(n5249), .B1(n2727), .B2(n2611), .ZN(n3969)
         );
  inv0d0 U4297 ( .I(\storage[7][7] ), .ZN(n2699) );
  aoi22d1 U4298 ( .A1(n2612), .A2(n3071), .B1(n2699), .B2(n2611), .ZN(n3968)
         );
  nr03d1 U4299 ( .A1(n2616), .A2(n2615), .A3(n2637), .ZN(n2617) );
  buffd1 U4300 ( .I(n2617), .Z(n2619) );
  aoim22d1 U4301 ( .A1(n2617), .A2(n266), .B1(\storage[6][0] ), .B2(n2619), 
        .Z(n3967) );
  inv0d0 U4302 ( .I(\storage[6][1] ), .ZN(n2824) );
  inv0d0 U4303 ( .I(n2619), .ZN(n2618) );
  aoi22d1 U4304 ( .A1(n2617), .A2(n4862), .B1(n2824), .B2(n2618), .ZN(n3966)
         );
  aoim22d1 U4305 ( .A1(n2617), .A2(n5004), .B1(\storage[6][2] ), .B2(n2619), 
        .Z(n3965) );
  aoim22d1 U4306 ( .A1(n2617), .A2(n5006), .B1(\storage[6][3] ), .B2(n2619), 
        .Z(n3964) );
  aoim22d1 U4307 ( .A1(n2617), .A2(n5008), .B1(\storage[6][4] ), .B2(n2619), 
        .Z(n3963) );
  aoim22d1 U4308 ( .A1(n2617), .A2(n5248), .B1(\storage[6][5] ), .B2(n2619), 
        .Z(n3962) );
  inv0d0 U4309 ( .I(\storage[6][6] ), .ZN(n2737) );
  aoi22d1 U4310 ( .A1(n2617), .A2(n2641), .B1(n2737), .B2(n2618), .ZN(n3961)
         );
  inv0d0 U4311 ( .I(\storage[6][7] ), .ZN(n2712) );
  aoi22d1 U4312 ( .A1(n2619), .A2(n3071), .B1(n2712), .B2(n2618), .ZN(n3960)
         );
  nr02d1 U4313 ( .A1(n2624), .A2(n2633), .ZN(n2623) );
  inv0d0 U4314 ( .I(\storage[5][0] ), .ZN(n2679) );
  inv0d0 U4315 ( .I(n2623), .ZN(n2622) );
  aoi22d1 U4316 ( .A1(n2623), .A2(n5290), .B1(n2679), .B2(n2622), .ZN(n3959)
         );
  inv0d0 U4317 ( .I(\storage[5][1] ), .ZN(n2815) );
  aoi22d1 U4318 ( .A1(n2623), .A2(n5294), .B1(n2815), .B2(n2622), .ZN(n3958)
         );
  aoim22d1 U4319 ( .A1(n2623), .A2(n5004), .B1(\storage[5][2] ), .B2(n2623), 
        .Z(n3957) );
  aoim22d1 U4320 ( .A1(n2623), .A2(n5006), .B1(\storage[5][3] ), .B2(n2623), 
        .Z(n3956) );
  aoim22d1 U4321 ( .A1(n2623), .A2(n5008), .B1(\storage[5][4] ), .B2(n2623), 
        .Z(n3955) );
  inv0d0 U4322 ( .I(\storage[5][5] ), .ZN(n2748) );
  aoi22d1 U4323 ( .A1(n2623), .A2(n2640), .B1(n2748), .B2(n2622), .ZN(n3954)
         );
  inv0d0 U4324 ( .I(\storage[5][6] ), .ZN(n2724) );
  aoi22d1 U4325 ( .A1(n2623), .A2(n5012), .B1(n2724), .B2(n2622), .ZN(n3953)
         );
  inv0d0 U4326 ( .I(\storage[5][7] ), .ZN(n2700) );
  aoi22d1 U4327 ( .A1(n2623), .A2(n3071), .B1(n2700), .B2(n2622), .ZN(n3952)
         );
  nr02d1 U4328 ( .A1(n2624), .A2(n2637), .ZN(n2627) );
  aoim22d1 U4329 ( .A1(n2627), .A2(n266), .B1(\storage[4][0] ), .B2(n2627), 
        .Z(n3951) );
  inv0d0 U4330 ( .I(\storage[4][1] ), .ZN(n2836) );
  inv0d0 U4331 ( .I(n2627), .ZN(n2626) );
  aoi22d1 U4332 ( .A1(n2627), .A2(n4862), .B1(n2836), .B2(n2626), .ZN(n3950)
         );
  aoim22d1 U4333 ( .A1(n2627), .A2(n5004), .B1(\storage[4][2] ), .B2(n2627), 
        .Z(n3949) );
  aoim22d1 U4334 ( .A1(n2627), .A2(n2625), .B1(\storage[4][3] ), .B2(n2627), 
        .Z(n3948) );
  aoim22d1 U4335 ( .A1(n2627), .A2(n4866), .B1(\storage[4][4] ), .B2(n2627), 
        .Z(n3947) );
  aoim22d1 U4336 ( .A1(n2627), .A2(n5010), .B1(\storage[4][5] ), .B2(n2627), 
        .Z(n3946) );
  inv0d0 U4337 ( .I(\storage[4][6] ), .ZN(n2734) );
  aoi22d1 U4338 ( .A1(n2627), .A2(n2641), .B1(n2734), .B2(n2626), .ZN(n3945)
         );
  inv0d0 U4339 ( .I(\storage[4][7] ), .ZN(n2711) );
  aoi22d1 U4340 ( .A1(n2627), .A2(n3071), .B1(n2711), .B2(n2626), .ZN(n3944)
         );
  nr02d1 U4341 ( .A1(n2630), .A2(n2633), .ZN(n2629) );
  inv0d0 U4342 ( .I(\storage[3][0] ), .ZN(n2675) );
  inv0d0 U4343 ( .I(n2629), .ZN(n2628) );
  aoi22d1 U4344 ( .A1(n2629), .A2(n4808), .B1(n2675), .B2(n2628), .ZN(n3943)
         );
  inv0d0 U4345 ( .I(\storage[3][1] ), .ZN(n2813) );
  aoi22d1 U4346 ( .A1(n2629), .A2(n4862), .B1(n2813), .B2(n2628), .ZN(n3942)
         );
  aoim22d1 U4347 ( .A1(n2629), .A2(n5245), .B1(\storage[3][2] ), .B2(n2629), 
        .Z(n3941) );
  aoim22d1 U4348 ( .A1(n2629), .A2(n5246), .B1(\storage[3][3] ), .B2(n2629), 
        .Z(n3940) );
  aoim22d1 U4349 ( .A1(n2629), .A2(n5247), .B1(\storage[3][4] ), .B2(n2629), 
        .Z(n3939) );
  inv0d0 U4350 ( .I(\storage[3][5] ), .ZN(n2753) );
  aoi22d1 U4351 ( .A1(n2629), .A2(n5010), .B1(n2753), .B2(n2628), .ZN(n3938)
         );
  inv0d0 U4352 ( .I(\storage[3][6] ), .ZN(n2729) );
  aoi22d1 U4353 ( .A1(n2629), .A2(n5249), .B1(n2729), .B2(n2628), .ZN(n3937)
         );
  inv0d0 U4354 ( .I(\storage[3][7] ), .ZN(n2698) );
  aoi22d1 U4355 ( .A1(n2629), .A2(n3071), .B1(n2698), .B2(n2628), .ZN(n3936)
         );
  nr02d1 U4356 ( .A1(n2630), .A2(n2637), .ZN(n2632) );
  aoim22d1 U4357 ( .A1(n2632), .A2(n4808), .B1(\storage[2][0] ), .B2(n2632), 
        .Z(n3935) );
  inv0d0 U4358 ( .I(\storage[2][1] ), .ZN(n2832) );
  inv0d0 U4359 ( .I(n2632), .ZN(n2631) );
  aoi22d1 U4360 ( .A1(n2632), .A2(n4862), .B1(n2832), .B2(n2631), .ZN(n3934)
         );
  aoim22d1 U4361 ( .A1(n2632), .A2(n5004), .B1(\storage[2][2] ), .B2(n2632), 
        .Z(n3933) );
  aoim22d1 U4362 ( .A1(n2632), .A2(n5246), .B1(\storage[2][3] ), .B2(n2632), 
        .Z(n3932) );
  aoim22d1 U4363 ( .A1(n2632), .A2(n5247), .B1(\storage[2][4] ), .B2(n2632), 
        .Z(n3931) );
  aoim22d1 U4364 ( .A1(n2632), .A2(n5010), .B1(\storage[2][5] ), .B2(n2632), 
        .Z(n3930) );
  inv0d0 U4365 ( .I(\storage[2][6] ), .ZN(n2736) );
  aoi22d1 U4366 ( .A1(n2632), .A2(n5249), .B1(n2736), .B2(n2631), .ZN(n3929)
         );
  inv0d0 U4367 ( .I(\storage[2][7] ), .ZN(n2713) );
  aoi22d1 U4368 ( .A1(n2632), .A2(n5251), .B1(n2713), .B2(n2631), .ZN(n3928)
         );
  nr02d1 U4369 ( .A1(n2638), .A2(n2633), .ZN(n2636) );
  inv0d0 U4370 ( .I(\storage[1][0] ), .ZN(n2678) );
  inv0d0 U4371 ( .I(n2636), .ZN(n2634) );
  aoi22d1 U4372 ( .A1(n2636), .A2(n5290), .B1(n2678), .B2(n2634), .ZN(n3927)
         );
  inv0d0 U4373 ( .I(\storage[1][1] ), .ZN(n2811) );
  aoi22d1 U4374 ( .A1(n2636), .A2(n5294), .B1(n2811), .B2(n2634), .ZN(n3926)
         );
  aoim22d1 U4375 ( .A1(n2636), .A2(n5245), .B1(\storage[1][2] ), .B2(n2636), 
        .Z(n3925) );
  aoim22d1 U4376 ( .A1(n2636), .A2(n5246), .B1(\storage[1][3] ), .B2(n2636), 
        .Z(n3924) );
  aoim22d1 U4377 ( .A1(n2636), .A2(n5247), .B1(\storage[1][4] ), .B2(n2636), 
        .Z(n3923) );
  inv0d0 U4378 ( .I(\storage[1][5] ), .ZN(n2752) );
  aoi22d1 U4379 ( .A1(n2636), .A2(n2640), .B1(n2752), .B2(n2634), .ZN(n3922)
         );
  inv0d0 U4380 ( .I(\storage[1][6] ), .ZN(n2728) );
  aoi22d1 U4381 ( .A1(n2636), .A2(n5012), .B1(n2728), .B2(n2634), .ZN(n3921)
         );
  inv0d0 U4382 ( .I(\storage[1][7] ), .ZN(n2696) );
  aoi22d1 U4383 ( .A1(n2636), .A2(n2635), .B1(n2696), .B2(n2634), .ZN(n3920)
         );
  nr02d1 U4384 ( .A1(n2638), .A2(n2637), .ZN(n2643) );
  aoim22d1 U4385 ( .A1(n2643), .A2(n266), .B1(\storage[0][0] ), .B2(n2643), 
        .Z(n3919) );
  inv0d0 U4386 ( .I(\storage[0][1] ), .ZN(n2828) );
  inv0d0 U4387 ( .I(n2643), .ZN(n2642) );
  aoi22d1 U4388 ( .A1(n2643), .A2(n2639), .B1(n2828), .B2(n2642), .ZN(n3918)
         );
  aoim22d1 U4389 ( .A1(n2643), .A2(n5004), .B1(\storage[0][2] ), .B2(n2643), 
        .Z(n3917) );
  aoim22d1 U4390 ( .A1(n2643), .A2(n5246), .B1(\storage[0][3] ), .B2(n2643), 
        .Z(n3916) );
  aoim22d1 U4391 ( .A1(n2643), .A2(n5247), .B1(\storage[0][4] ), .B2(n2643), 
        .Z(n3915) );
  aoim22d1 U4392 ( .A1(n2643), .A2(n2640), .B1(\storage[0][5] ), .B2(n2643), 
        .Z(n3914) );
  inv0d0 U4393 ( .I(\storage[0][6] ), .ZN(n2738) );
  aoi22d1 U4394 ( .A1(n2643), .A2(n2641), .B1(n2738), .B2(n2642), .ZN(n3913)
         );
  inv0d0 U4395 ( .I(\storage[0][7] ), .ZN(n2709) );
  aoi22d1 U4396 ( .A1(n2643), .A2(n5251), .B1(n2709), .B2(n2642), .ZN(n3912)
         );
  inv0d0 U4397 ( .I(n2644), .ZN(n2645) );
  aoi21d1 U4398 ( .B1(n2646), .B2(n2645), .A(n5111), .ZN(n3911) );
  oai21d1 U4399 ( .B1(n2655), .B2(n4575), .A(n5319), .ZN(n2651) );
  nd02d0 U4400 ( .A1(n2648), .A2(n2647), .ZN(n2652) );
  inv0d0 U4401 ( .I(csrbank11_ev_enable0_w[0]), .ZN(n2649) );
  aoi22d1 U4402 ( .A1(n5000), .A2(n2651), .B1(n2652), .B2(n2649), .ZN(n3910)
         );
  inv0d0 U4403 ( .I(csrbank11_ev_enable0_w[1]), .ZN(n2650) );
  oai22d1 U4404 ( .A1(n2653), .A2(n2652), .B1(n2651), .B2(n2650), .ZN(n3909)
         );
  inv0d0 U4405 ( .I(N5711), .ZN(n2659) );
  inv0d0 U4406 ( .I(uart_pending_r[0]), .ZN(n2656) );
  oai21d1 U4407 ( .B1(n2655), .B2(n2654), .A(n5319), .ZN(n2658) );
  oai22d1 U4408 ( .A1(n4808), .A2(n2659), .B1(n2656), .B2(n2658), .ZN(n3908)
         );
  inv0d0 U4409 ( .I(uart_pending_r[1]), .ZN(n2657) );
  oai22d1 U4410 ( .A1(n4862), .A2(n2659), .B1(n2658), .B2(n2657), .ZN(n3907)
         );
  nd02d0 U4411 ( .A1(uart_pending_status[1]), .A2(n2660), .ZN(n2661) );
  oan211d1 U4412 ( .C1(uart_rx_trigger_d), .C2(n2662), .B(n2661), .A(n5492), 
        .ZN(n3906) );
  oaim21d1 U4413 ( .B1(uart_pending_r[0]), .B2(uart_pending_re), .A(
        uart_pending_status[0]), .ZN(n2663) );
  oan211d1 U4414 ( .C1(n2664), .C2(uart_tx_trigger_d), .B(n2663), .A(n2516), 
        .ZN(n3905) );
  aoi211d1 U4415 ( .C1(n2666), .C2(n2848), .A(n4878), .B(n2665), .ZN(n3904) );
  inv0d0 U4416 ( .I(uart_phy_tx_tick), .ZN(n2867) );
  inv0d0 U4417 ( .I(uart_phy_tx_count[0]), .ZN(n2667) );
  aoi221d1 U4418 ( .B1(uart_phy_tx_tick), .B2(uart_phy_tx_count[0]), .C1(n2867), .C2(n2667), .A(n2848), .ZN(n3903) );
  inv0d0 U4419 ( .I(uart_phy_tx_count[1]), .ZN(n2668) );
  aoi211d1 U4420 ( .C1(n2669), .C2(n2668), .A(n2673), .B(n2848), .ZN(n3902) );
  inv0d0 U4421 ( .I(n2673), .ZN(n2670) );
  aoi221d1 U4422 ( .B1(uart_phy_tx_count[2]), .B2(n2673), .C1(n2671), .C2(
        n2670), .A(n2848), .ZN(n3901) );
  aon211d1 U4423 ( .C1(uart_phy_tx_count[2]), .C2(n2673), .B(
        uart_phy_tx_count[3]), .A(n2868), .ZN(n2672) );
  aoi31d1 U4424 ( .B1(uart_phy_tx_count[3]), .B2(uart_phy_tx_count[2]), .B3(
        n2673), .A(n2672), .ZN(n3900) );
  nr03d1 U4425 ( .A1(uart_tx_fifo_rdport_adr[3]), .A2(n2674), .A3(n2677), .ZN(
        n2795) );
  nr03d1 U4426 ( .A1(uart_tx_fifo_rdport_adr[1]), .A2(n2677), .A3(n2680), .ZN(
        n2797) );
  aoi22d1 U4427 ( .A1(\storage[7][0] ), .A2(n2795), .B1(\storage[13][0] ), 
        .B2(n2797), .ZN(n2693) );
  nr03d1 U4428 ( .A1(uart_tx_fifo_rdport_adr[2]), .A2(n2674), .A3(n2680), .ZN(
        n2799) );
  inv0d0 U4429 ( .I(n2799), .ZN(n2825) );
  nr03d0 U4430 ( .A1(uart_tx_fifo_rdport_adr[2]), .A2(
        uart_tx_fifo_rdport_adr[3]), .A3(n2674), .ZN(n2794) );
  inv0d0 U4431 ( .I(n2794), .ZN(n2831) );
  oai22d1 U4432 ( .A1(n2676), .A2(n2825), .B1(n2675), .B2(n2831), .ZN(n2685)
         );
  nr03d0 U4433 ( .A1(uart_tx_fifo_rdport_adr[1]), .A2(
        uart_tx_fifo_rdport_adr[3]), .A3(n2677), .ZN(n2800) );
  inv0d0 U4434 ( .I(n2800), .ZN(n2835) );
  nr03d0 U4435 ( .A1(uart_tx_fifo_rdport_adr[2]), .A2(
        uart_tx_fifo_rdport_adr[1]), .A3(uart_tx_fifo_rdport_adr[3]), .ZN(
        n2798) );
  inv0d0 U4436 ( .I(n2798), .ZN(n2827) );
  oai22d1 U4437 ( .A1(n2679), .A2(n2835), .B1(n2678), .B2(n2827), .ZN(n2684)
         );
  inv0d0 U4438 ( .I(n2801), .ZN(n2833) );
  nr03d0 U4439 ( .A1(uart_tx_fifo_rdport_adr[2]), .A2(
        uart_tx_fifo_rdport_adr[1]), .A3(n2680), .ZN(n2796) );
  inv0d0 U4440 ( .I(n2796), .ZN(n2829) );
  oai22d1 U4441 ( .A1(n2682), .A2(n2833), .B1(n2681), .B2(n2829), .ZN(n2683)
         );
  inv0d0 U4442 ( .I(n2767), .ZN(n2847) );
  nr02d0 U4443 ( .A1(uart_tx_fifo_rdport_adr[0]), .A2(n2809), .ZN(n2706) );
  aoi22d1 U4444 ( .A1(\storage[14][0] ), .A2(n2801), .B1(\storage[10][0] ), 
        .B2(n2799), .ZN(n2689) );
  aoi22d1 U4445 ( .A1(\storage[12][0] ), .A2(n2797), .B1(\storage[0][0] ), 
        .B2(n2798), .ZN(n2688) );
  aoi22d1 U4446 ( .A1(\storage[4][0] ), .A2(n2800), .B1(\storage[2][0] ), .B2(
        n2794), .ZN(n2687) );
  aoi22d1 U4447 ( .A1(\storage[8][0] ), .A2(n2796), .B1(\storage[6][0] ), .B2(
        n2795), .ZN(n2686) );
  aoi22d1 U4448 ( .A1(n2706), .A2(n2690), .B1(
        uart_tx_fifo_fifo_out_payload_data[0]), .B2(n2809), .ZN(n2691) );
  aon211d1 U4449 ( .C1(n2693), .C2(n2692), .B(n2847), .A(n2691), .ZN(n3899) );
  oai22d1 U4450 ( .A1(n2695), .A2(n2833), .B1(n2694), .B2(n2825), .ZN(n2705)
         );
  oai22d1 U4451 ( .A1(n2697), .A2(n2829), .B1(n2696), .B2(n2827), .ZN(n2704)
         );
  inv0d0 U4452 ( .I(n2795), .ZN(n2823) );
  oai22d1 U4453 ( .A1(n2699), .A2(n2823), .B1(n2698), .B2(n2831), .ZN(n2703)
         );
  inv0d0 U4454 ( .I(n2797), .ZN(n2837) );
  oai22d1 U4455 ( .A1(n2701), .A2(n2837), .B1(n2700), .B2(n2835), .ZN(n2702)
         );
  nr04d0 U4456 ( .A1(n2705), .A2(n2704), .A3(n2703), .A4(n2702), .ZN(n2721) );
  inv0d0 U4457 ( .I(uart_tx_fifo_fifo_out_payload_data[7]), .ZN(n2720) );
  inv0d0 U4458 ( .I(n2706), .ZN(n2844) );
  oai22d1 U4459 ( .A1(n2708), .A2(n2837), .B1(n2707), .B2(n2825), .ZN(n2718)
         );
  oai22d1 U4460 ( .A1(n2710), .A2(n2829), .B1(n2709), .B2(n2827), .ZN(n2717)
         );
  oai22d1 U4461 ( .A1(n2712), .A2(n2823), .B1(n2711), .B2(n2835), .ZN(n2716)
         );
  oai22d1 U4462 ( .A1(n2714), .A2(n2833), .B1(n2713), .B2(n2831), .ZN(n2715)
         );
  nr04d0 U4463 ( .A1(n2718), .A2(n2717), .A3(n2716), .A4(n2715), .ZN(n2719) );
  oai222d1 U4464 ( .A1(n2847), .A2(n2721), .B1(n2720), .B2(n2845), .C1(n2844), 
        .C2(n2719), .ZN(n3898) );
  oai22d1 U4465 ( .A1(n2723), .A2(n2833), .B1(n2722), .B2(n2837), .ZN(n2733)
         );
  oai22d1 U4466 ( .A1(n2725), .A2(n2825), .B1(n2724), .B2(n2835), .ZN(n2732)
         );
  oai22d1 U4467 ( .A1(n2727), .A2(n2823), .B1(n2726), .B2(n2829), .ZN(n2731)
         );
  oai22d1 U4468 ( .A1(n2729), .A2(n2831), .B1(n2728), .B2(n2827), .ZN(n2730)
         );
  nr04d0 U4469 ( .A1(n2733), .A2(n2732), .A3(n2731), .A4(n2730), .ZN(n2747) );
  inv0d0 U4470 ( .I(uart_tx_fifo_fifo_out_payload_data[6]), .ZN(n2861) );
  oai22d1 U4471 ( .A1(n2735), .A2(n2833), .B1(n2734), .B2(n2835), .ZN(n2745)
         );
  oai22d1 U4472 ( .A1(n2737), .A2(n2823), .B1(n2736), .B2(n2831), .ZN(n2744)
         );
  oai22d1 U4473 ( .A1(n2739), .A2(n2837), .B1(n2738), .B2(n2827), .ZN(n2743)
         );
  oai22d1 U4474 ( .A1(n2741), .A2(n2825), .B1(n2740), .B2(n2829), .ZN(n2742)
         );
  nr04d0 U4475 ( .A1(n2745), .A2(n2744), .A3(n2743), .A4(n2742), .ZN(n2746) );
  oai222d1 U4476 ( .A1(n2847), .A2(n2747), .B1(n2861), .B2(n2845), .C1(n2844), 
        .C2(n2746), .ZN(n3897) );
  oai22d1 U4477 ( .A1(n2749), .A2(n2833), .B1(n2748), .B2(n2835), .ZN(n2759)
         );
  oai22d1 U4478 ( .A1(n2751), .A2(n2823), .B1(n2750), .B2(n2825), .ZN(n2758)
         );
  oai22d1 U4479 ( .A1(n2753), .A2(n2831), .B1(n2752), .B2(n2827), .ZN(n2757)
         );
  oai22d1 U4480 ( .A1(n2755), .A2(n2837), .B1(n2754), .B2(n2829), .ZN(n2756)
         );
  aoi22d1 U4481 ( .A1(\storage[14][5] ), .A2(n2801), .B1(\storage[4][5] ), 
        .B2(n2800), .ZN(n2763) );
  aoi22d1 U4482 ( .A1(\storage[12][5] ), .A2(n2797), .B1(\storage[8][5] ), 
        .B2(n2796), .ZN(n2762) );
  aoi22d1 U4483 ( .A1(\storage[10][5] ), .A2(n2799), .B1(\storage[2][5] ), 
        .B2(n2794), .ZN(n2761) );
  aoi22d1 U4484 ( .A1(\storage[6][5] ), .A2(n2795), .B1(\storage[0][5] ), .B2(
        n2798), .ZN(n2760) );
  oai22d1 U4485 ( .A1(n2845), .A2(uart_tx_fifo_fifo_out_payload_data[5]), .B1(
        n2764), .B2(n2844), .ZN(n2765) );
  aoi21d1 U4486 ( .B1(n2767), .B2(n2766), .A(n2765), .ZN(n3896) );
  aoi22d1 U4487 ( .A1(\storage[11][4] ), .A2(n2799), .B1(\storage[9][4] ), 
        .B2(n2796), .ZN(n2771) );
  aoi22d1 U4488 ( .A1(\storage[13][4] ), .A2(n2797), .B1(\storage[5][4] ), 
        .B2(n2800), .ZN(n2770) );
  aoi22d1 U4489 ( .A1(\storage[15][4] ), .A2(n2801), .B1(\storage[1][4] ), 
        .B2(n2798), .ZN(n2769) );
  aoi22d1 U4490 ( .A1(\storage[7][4] ), .A2(n2795), .B1(\storage[3][4] ), .B2(
        n2794), .ZN(n2768) );
  aoi22d1 U4491 ( .A1(\storage[12][4] ), .A2(n2797), .B1(\storage[8][4] ), 
        .B2(n2796), .ZN(n2775) );
  aoi22d1 U4492 ( .A1(\storage[14][4] ), .A2(n2801), .B1(\storage[2][4] ), 
        .B2(n2794), .ZN(n2774) );
  aoi22d1 U4493 ( .A1(\storage[10][4] ), .A2(n2799), .B1(\storage[0][4] ), 
        .B2(n2798), .ZN(n2773) );
  aoi22d1 U4494 ( .A1(\storage[6][4] ), .A2(n2795), .B1(\storage[4][4] ), .B2(
        n2800), .ZN(n2772) );
  aoi22d1 U4495 ( .A1(uart_tx_fifo_rdport_adr[0]), .A2(n2777), .B1(n2776), 
        .B2(n2806), .ZN(n2778) );
  inv0d0 U4496 ( .I(uart_tx_fifo_fifo_out_payload_data[4]), .ZN(n2857) );
  aoi22d1 U4497 ( .A1(n2845), .A2(n2778), .B1(n2857), .B2(n2809), .ZN(n3895)
         );
  aoi22d1 U4498 ( .A1(\storage[13][3] ), .A2(n2797), .B1(\storage[3][3] ), 
        .B2(n2794), .ZN(n2782) );
  aoi22d1 U4499 ( .A1(\storage[7][3] ), .A2(n2795), .B1(\storage[5][3] ), .B2(
        n2800), .ZN(n2781) );
  aoi22d1 U4500 ( .A1(\storage[15][3] ), .A2(n2801), .B1(\storage[9][3] ), 
        .B2(n2796), .ZN(n2780) );
  aoi22d1 U4501 ( .A1(\storage[11][3] ), .A2(n2799), .B1(\storage[1][3] ), 
        .B2(n2798), .ZN(n2779) );
  aoi22d1 U4502 ( .A1(\storage[14][3] ), .A2(n2801), .B1(\storage[4][3] ), 
        .B2(n2800), .ZN(n2786) );
  aoi22d1 U4503 ( .A1(\storage[8][3] ), .A2(n2796), .B1(\storage[2][3] ), .B2(
        n2794), .ZN(n2785) );
  aoi22d1 U4504 ( .A1(\storage[12][3] ), .A2(n2797), .B1(\storage[10][3] ), 
        .B2(n2799), .ZN(n2784) );
  aoi22d1 U4505 ( .A1(\storage[6][3] ), .A2(n2795), .B1(\storage[0][3] ), .B2(
        n2798), .ZN(n2783) );
  aoi22d1 U4506 ( .A1(uart_tx_fifo_rdport_adr[0]), .A2(n2788), .B1(n2787), 
        .B2(n2806), .ZN(n2789) );
  inv0d0 U4507 ( .I(uart_tx_fifo_fifo_out_payload_data[3]), .ZN(n2855) );
  aoi22d1 U4508 ( .A1(n2845), .A2(n2789), .B1(n2855), .B2(n2809), .ZN(n3894)
         );
  aoi22d1 U4509 ( .A1(\storage[13][2] ), .A2(n2797), .B1(\storage[5][2] ), 
        .B2(n2800), .ZN(n2793) );
  aoi22d1 U4510 ( .A1(\storage[7][2] ), .A2(n2795), .B1(\storage[3][2] ), .B2(
        n2794), .ZN(n2792) );
  aoi22d1 U4511 ( .A1(\storage[11][2] ), .A2(n2799), .B1(\storage[9][2] ), 
        .B2(n2796), .ZN(n2791) );
  aoi22d1 U4512 ( .A1(\storage[15][2] ), .A2(n2801), .B1(\storage[1][2] ), 
        .B2(n2798), .ZN(n2790) );
  aoi22d1 U4513 ( .A1(\storage[6][2] ), .A2(n2795), .B1(\storage[2][2] ), .B2(
        n2794), .ZN(n2805) );
  aoi22d1 U4514 ( .A1(\storage[12][2] ), .A2(n2797), .B1(\storage[8][2] ), 
        .B2(n2796), .ZN(n2804) );
  aoi22d1 U4515 ( .A1(\storage[10][2] ), .A2(n2799), .B1(\storage[0][2] ), 
        .B2(n2798), .ZN(n2803) );
  aoi22d1 U4516 ( .A1(\storage[14][2] ), .A2(n2801), .B1(\storage[4][2] ), 
        .B2(n2800), .ZN(n2802) );
  aoi22d1 U4517 ( .A1(uart_tx_fifo_rdport_adr[0]), .A2(n2808), .B1(n2807), 
        .B2(n2806), .ZN(n2810) );
  inv0d0 U4518 ( .I(uart_tx_fifo_fifo_out_payload_data[2]), .ZN(n2853) );
  aoi22d1 U4519 ( .A1(n2845), .A2(n2810), .B1(n2853), .B2(n2809), .ZN(n3893)
         );
  oai22d1 U4520 ( .A1(n2812), .A2(n2825), .B1(n2811), .B2(n2827), .ZN(n2822)
         );
  oai22d1 U4521 ( .A1(n2814), .A2(n2833), .B1(n2813), .B2(n2831), .ZN(n2821)
         );
  oai22d1 U4522 ( .A1(n2816), .A2(n2829), .B1(n2815), .B2(n2835), .ZN(n2820)
         );
  oai22d1 U4523 ( .A1(n2818), .A2(n2823), .B1(n2817), .B2(n2837), .ZN(n2819)
         );
  nr04d0 U4524 ( .A1(n2822), .A2(n2821), .A3(n2820), .A4(n2819), .ZN(n2846) );
  inv0d0 U4525 ( .I(uart_tx_fifo_fifo_out_payload_data[1]), .ZN(n2851) );
  oai22d1 U4526 ( .A1(n2826), .A2(n2825), .B1(n2824), .B2(n2823), .ZN(n2842)
         );
  oai22d1 U4527 ( .A1(n2830), .A2(n2829), .B1(n2828), .B2(n2827), .ZN(n2841)
         );
  oai22d1 U4528 ( .A1(n2834), .A2(n2833), .B1(n2832), .B2(n2831), .ZN(n2840)
         );
  oai22d1 U4529 ( .A1(n2838), .A2(n2837), .B1(n2836), .B2(n2835), .ZN(n2839)
         );
  oai222d1 U4530 ( .A1(n2847), .A2(n2846), .B1(n2851), .B2(n2845), .C1(n2844), 
        .C2(n2843), .ZN(n3892) );
  inv0d0 U4531 ( .I(uart_phy_tx_data[1]), .ZN(n2850) );
  nd02d0 U4532 ( .A1(rs232phy_rs232phytx_state), .A2(uart_phy_tx_tick), .ZN(
        n2870) );
  nd02d0 U4533 ( .A1(uart_phy_tx_sink_valid), .A2(n2848), .ZN(n2864) );
  inv0d0 U4534 ( .I(uart_tx_fifo_fifo_out_payload_data[0]), .ZN(n2849) );
  nd02d0 U4535 ( .A1(n2870), .A2(n2864), .ZN(n2863) );
  inv0d0 U4536 ( .I(uart_phy_tx_data[0]), .ZN(n2871) );
  oai222d1 U4537 ( .A1(n2850), .A2(n2870), .B1(n2864), .B2(n2849), .C1(n2863), 
        .C2(n2871), .ZN(n3891) );
  inv0d0 U4538 ( .I(uart_phy_tx_data[2]), .ZN(n2852) );
  oai222d1 U4539 ( .A1(n2852), .A2(n2870), .B1(n2864), .B2(n2851), .C1(n2850), 
        .C2(n2863), .ZN(n3890) );
  inv0d0 U4540 ( .I(uart_phy_tx_data[3]), .ZN(n2854) );
  oai222d1 U4541 ( .A1(n2854), .A2(n2870), .B1(n2864), .B2(n2853), .C1(n2852), 
        .C2(n2863), .ZN(n3889) );
  inv0d0 U4542 ( .I(uart_phy_tx_data[4]), .ZN(n2856) );
  oai222d1 U4543 ( .A1(n2856), .A2(n2870), .B1(n2864), .B2(n2855), .C1(n2854), 
        .C2(n2863), .ZN(n3888) );
  inv0d0 U4544 ( .I(uart_phy_tx_data[5]), .ZN(n2858) );
  oai222d1 U4545 ( .A1(n2858), .A2(n2870), .B1(n2864), .B2(n2857), .C1(n2856), 
        .C2(n2863), .ZN(n3887) );
  inv0d0 U4546 ( .I(uart_phy_tx_data[6]), .ZN(n2860) );
  inv0d0 U4547 ( .I(uart_tx_fifo_fifo_out_payload_data[5]), .ZN(n2859) );
  oai222d1 U4548 ( .A1(n2860), .A2(n2870), .B1(n2864), .B2(n2859), .C1(n2858), 
        .C2(n2863), .ZN(n3886) );
  inv0d0 U4549 ( .I(uart_phy_tx_data[7]), .ZN(n2862) );
  oai222d1 U4550 ( .A1(n2862), .A2(n2870), .B1(n2864), .B2(n2861), .C1(n2860), 
        .C2(n2863), .ZN(n3885) );
  oai22d1 U4551 ( .A1(n2864), .A2(uart_tx_fifo_fifo_out_payload_data[7]), .B1(
        n2863), .B2(uart_phy_tx_data[7]), .ZN(n2865) );
  inv0d0 U4552 ( .I(n2865), .ZN(n3884) );
  oai21d1 U4553 ( .B1(uart_phy_tx_sink_valid), .B2(n2868), .A(n5319), .ZN(
        n2866) );
  aoi31d1 U4554 ( .B1(n2868), .B2(sys_uart_tx), .B3(n2867), .A(n2866), .ZN(
        n2869) );
  oai21d1 U4555 ( .B1(n2871), .B2(n2870), .A(n2869), .ZN(n3883) );
  ora211d1 U4556 ( .C1(dbg_uart_rx_tick), .C2(dbg_uart_rx_count[0]), .A(n2872), 
        .B(uartwishbonebridge_rs232phyrx_state), .Z(n3881) );
  nd02d0 U4557 ( .A1(n2873), .A2(dbg_uart_rx_count[2]), .ZN(n2875) );
  inv0d0 U4558 ( .I(n2875), .ZN(n2877) );
  aoim211d1 U4559 ( .C1(n2873), .C2(dbg_uart_rx_count[2]), .A(n2877), .B(n2874), .ZN(n3879) );
  aoi221d1 U4560 ( .B1(dbg_uart_rx_count[3]), .B2(n2877), .C1(n2876), .C2(
        n2875), .A(n2874), .ZN(n3878) );
  nd02d0 U4561 ( .A1(dbg_uart_rx_tick), .A2(
        uartwishbonebridge_rs232phyrx_state), .ZN(n2878) );
  inv0d0 U4562 ( .I(n2878), .ZN(n2880) );
  inv0d0 U4563 ( .I(dbg_uart_rx_data[1]), .ZN(n5970) );
  inv0d0 U4564 ( .I(dbg_uart_rx_data[0]), .ZN(n5969) );
  aoi22d1 U4565 ( .A1(n2880), .A2(n5970), .B1(n5969), .B2(n2878), .ZN(n3877)
         );
  inv0d0 U4566 ( .I(dbg_uart_rx_data[2]), .ZN(n5971) );
  aoi22d1 U4567 ( .A1(n2880), .A2(n5971), .B1(n5970), .B2(n2878), .ZN(n3876)
         );
  inv0d0 U4568 ( .I(dbg_uart_rx_data[3]), .ZN(n5972) );
  aoi22d1 U4569 ( .A1(n2880), .A2(n5972), .B1(n5971), .B2(n2878), .ZN(n3875)
         );
  inv0d0 U4570 ( .I(dbg_uart_rx_data[4]), .ZN(n5973) );
  aoi22d1 U4571 ( .A1(n2880), .A2(n5973), .B1(n5972), .B2(n2878), .ZN(n3874)
         );
  inv0d0 U4572 ( .I(dbg_uart_rx_data[5]), .ZN(n5974) );
  aoi22d1 U4573 ( .A1(n2880), .A2(n5974), .B1(n5973), .B2(n2878), .ZN(n3873)
         );
  inv0d0 U4574 ( .I(dbg_uart_rx_data[6]), .ZN(n5975) );
  aoi22d1 U4575 ( .A1(n2880), .A2(n5975), .B1(n5974), .B2(n2878), .ZN(n3872)
         );
  inv0d0 U4576 ( .I(dbg_uart_rx_data[7]), .ZN(n5976) );
  aoi22d1 U4577 ( .A1(n2880), .A2(n5976), .B1(n5975), .B2(n2878), .ZN(n3871)
         );
  aoi22d1 U4578 ( .A1(n2880), .A2(n2879), .B1(n5976), .B2(n2878), .ZN(n3870)
         );
  inv0d0 U4579 ( .I(uart_phy_rx_tick), .ZN(n2882) );
  inv0d0 U4580 ( .I(uart_phy_rx_count[0]), .ZN(n2881) );
  oai21d1 U4581 ( .B1(n2882), .B2(n2881), .A(rs232phy_rs232phyrx_state), .ZN(
        n2883) );
  aoi21d1 U4582 ( .B1(n2882), .B2(n2881), .A(n2883), .ZN(n3868) );
  inv0d0 U4583 ( .I(uart_phy_rx_count[1]), .ZN(n2886) );
  aoi22d1 U4584 ( .A1(uart_phy_rx_count[1]), .A2(n2883), .B1(n2889), .B2(n2886), .ZN(n3867) );
  inv0d0 U4585 ( .I(uart_phy_rx_count[2]), .ZN(n2885) );
  nd02d0 U4586 ( .A1(uart_phy_rx_count[1]), .A2(uart_phy_rx_count[2]), .ZN(
        n2888) );
  inv0d0 U4587 ( .I(n2883), .ZN(n2884) );
  aoi21d1 U4588 ( .B1(rs232phy_rs232phyrx_state), .B2(n2888), .A(n2884), .ZN(
        n2887) );
  oan211d1 U4589 ( .C1(n2889), .C2(n2886), .B(n2885), .A(n2887), .ZN(n3866) );
  aoi222d1 U4590 ( .A1(n2890), .A2(n2889), .B1(n2890), .B2(n2888), .C1(
        uart_phy_rx_count[3]), .C2(n2887), .ZN(n3865) );
  inv0d1 U4591 ( .I(uart_phy_rx_data[0]), .ZN(n3047) );
  inv0d0 U4592 ( .I(n2893), .ZN(n2892) );
  aoi22d1 U4593 ( .A1(n2893), .A2(n3047), .B1(n2891), .B2(n2892), .ZN(n3864)
         );
  aoim22d1 U4594 ( .A1(n2893), .A2(n3048), .B1(\storage_1[15][1] ), .B2(n2893), 
        .Z(n3863) );
  aoim22d1 U4595 ( .A1(n2893), .A2(n3049), .B1(\storage_1[15][2] ), .B2(n2893), 
        .Z(n3862) );
  aoim22d1 U4596 ( .A1(n2893), .A2(n3050), .B1(\storage_1[15][3] ), .B2(n2893), 
        .Z(n3861) );
  inv0d0 U4597 ( .I(\storage_1[15][4] ), .ZN(n2972) );
  aoi22d1 U4598 ( .A1(n2893), .A2(n3051), .B1(n2972), .B2(n2892), .ZN(n3860)
         );
  aoim22d1 U4599 ( .A1(n2893), .A2(n3052), .B1(\storage_1[15][5] ), .B2(n2893), 
        .Z(n3859) );
  inv0d0 U4600 ( .I(\storage_1[15][6] ), .ZN(n3004) );
  aoi22d1 U4601 ( .A1(n2893), .A2(n3053), .B1(n3004), .B2(n2892), .ZN(n3858)
         );
  aoim22d1 U4602 ( .A1(n2893), .A2(n3055), .B1(\storage_1[15][7] ), .B2(n2893), 
        .Z(n3857) );
  nd03d0 U4603 ( .A1(uart_rx_fifo_produce[3]), .A2(n2915), .A3(n2913), .ZN(
        n2907) );
  nr02d1 U4604 ( .A1(n2916), .A2(n2907), .ZN(n2894) );
  aoim22d1 U4605 ( .A1(n2894), .A2(n3047), .B1(\storage_1[14][0] ), .B2(n2894), 
        .Z(n3856) );
  aoim22d1 U4606 ( .A1(n2894), .A2(n3048), .B1(\storage_1[14][1] ), .B2(n2894), 
        .Z(n3855) );
  aoim22d1 U4607 ( .A1(n2894), .A2(n3049), .B1(\storage_1[14][2] ), .B2(n2894), 
        .Z(n3854) );
  aoim22d1 U4608 ( .A1(n2894), .A2(n3050), .B1(\storage_1[14][3] ), .B2(n2894), 
        .Z(n3853) );
  aoim22d1 U4609 ( .A1(n2894), .A2(n3051), .B1(\storage_1[14][4] ), .B2(n2894), 
        .Z(n3852) );
  aoim22d1 U4610 ( .A1(n2894), .A2(n3052), .B1(\storage_1[14][5] ), .B2(n2894), 
        .Z(n3851) );
  aoim22d1 U4611 ( .A1(n2894), .A2(n3053), .B1(\storage_1[14][6] ), .B2(n2894), 
        .Z(n3850) );
  aoim22d1 U4612 ( .A1(n2894), .A2(n3055), .B1(\storage_1[14][7] ), .B2(n2894), 
        .Z(n3849) );
  nd02d0 U4613 ( .A1(uart_rx_fifo_produce[2]), .A2(n2901), .ZN(n2921) );
  nr02d1 U4614 ( .A1(n2903), .A2(n2921), .ZN(n2897) );
  inv0d0 U4615 ( .I(n2897), .ZN(n2896) );
  aoi22d1 U4616 ( .A1(n2897), .A2(n3047), .B1(n2895), .B2(n2896), .ZN(n3848)
         );
  aoim22d1 U4617 ( .A1(n2897), .A2(n3048), .B1(\storage_1[13][1] ), .B2(n2897), 
        .Z(n3847) );
  aoim22d1 U4618 ( .A1(n2897), .A2(n3049), .B1(\storage_1[13][2] ), .B2(n2897), 
        .Z(n3846) );
  aoim22d1 U4619 ( .A1(n2897), .A2(n3050), .B1(\storage_1[13][3] ), .B2(n2897), 
        .Z(n3845) );
  inv0d0 U4620 ( .I(\storage_1[13][4] ), .ZN(n2971) );
  aoi22d1 U4621 ( .A1(n2897), .A2(n3051), .B1(n2971), .B2(n2896), .ZN(n3844)
         );
  aoim22d1 U4622 ( .A1(n2897), .A2(n3052), .B1(\storage_1[13][5] ), .B2(n2897), 
        .Z(n3843) );
  inv0d0 U4623 ( .I(\storage_1[13][6] ), .ZN(n3008) );
  aoi22d1 U4624 ( .A1(n2897), .A2(n3053), .B1(n3008), .B2(n2896), .ZN(n3842)
         );
  aoim22d1 U4625 ( .A1(n2897), .A2(n3055), .B1(\storage_1[13][7] ), .B2(n2897), 
        .Z(n3841) );
  nr02d1 U4626 ( .A1(n2907), .A2(n2921), .ZN(n2898) );
  aoim22d1 U4627 ( .A1(n2898), .A2(n3047), .B1(\storage_1[12][0] ), .B2(n2898), 
        .Z(n3840) );
  aoim22d1 U4628 ( .A1(n2898), .A2(n3048), .B1(\storage_1[12][1] ), .B2(n2898), 
        .Z(n3839) );
  aoim22d1 U4629 ( .A1(n2898), .A2(n3049), .B1(\storage_1[12][2] ), .B2(n2898), 
        .Z(n3838) );
  aoim22d1 U4630 ( .A1(n2898), .A2(n3050), .B1(\storage_1[12][3] ), .B2(n2898), 
        .Z(n3837) );
  aoim22d1 U4631 ( .A1(n2898), .A2(n3051), .B1(\storage_1[12][4] ), .B2(n2898), 
        .Z(n3836) );
  aoim22d1 U4632 ( .A1(n2898), .A2(n3052), .B1(\storage_1[12][5] ), .B2(n2898), 
        .Z(n3835) );
  aoim22d1 U4633 ( .A1(n2898), .A2(n3053), .B1(\storage_1[12][6] ), .B2(n2898), 
        .Z(n3834) );
  aoim22d1 U4634 ( .A1(n2898), .A2(n3055), .B1(\storage_1[12][7] ), .B2(n2898), 
        .Z(n3833) );
  nd02d0 U4635 ( .A1(uart_rx_fifo_produce[1]), .A2(n2902), .ZN(n2924) );
  nr02d1 U4636 ( .A1(n2903), .A2(n2924), .ZN(n2899) );
  aoim22d1 U4637 ( .A1(n2899), .A2(n3047), .B1(\storage_1[11][0] ), .B2(n2899), 
        .Z(n3832) );
  aoim22d1 U4638 ( .A1(n2899), .A2(n3048), .B1(\storage_1[11][1] ), .B2(n2899), 
        .Z(n3831) );
  aoim22d1 U4639 ( .A1(n2899), .A2(n3049), .B1(\storage_1[11][2] ), .B2(n2899), 
        .Z(n3830) );
  aoim22d1 U4640 ( .A1(n2899), .A2(n3050), .B1(\storage_1[11][3] ), .B2(n2899), 
        .Z(n3829) );
  aoim22d1 U4641 ( .A1(n2899), .A2(n3051), .B1(\storage_1[11][4] ), .B2(n2899), 
        .Z(n3828) );
  aoim22d1 U4642 ( .A1(n2899), .A2(n3052), .B1(\storage_1[11][5] ), .B2(n2899), 
        .Z(n3827) );
  aoim22d1 U4643 ( .A1(n2899), .A2(n3053), .B1(\storage_1[11][6] ), .B2(n2899), 
        .Z(n3826) );
  aoim22d1 U4644 ( .A1(n2899), .A2(n3055), .B1(\storage_1[11][7] ), .B2(n2899), 
        .Z(n3825) );
  nr02d1 U4645 ( .A1(n2907), .A2(n2924), .ZN(n2900) );
  aoim22d1 U4646 ( .A1(n2900), .A2(n3047), .B1(\storage_1[10][0] ), .B2(n2900), 
        .Z(n3824) );
  aoim22d1 U4647 ( .A1(n2900), .A2(n3048), .B1(\storage_1[10][1] ), .B2(n2900), 
        .Z(n3823) );
  aoim22d1 U4648 ( .A1(n2900), .A2(n3049), .B1(\storage_1[10][2] ), .B2(n2900), 
        .Z(n3822) );
  aoim22d1 U4649 ( .A1(n2900), .A2(n3050), .B1(\storage_1[10][3] ), .B2(n2900), 
        .Z(n3821) );
  aoim22d1 U4650 ( .A1(n2900), .A2(n3051), .B1(\storage_1[10][4] ), .B2(n2900), 
        .Z(n3820) );
  aoim22d1 U4651 ( .A1(n2900), .A2(n3052), .B1(\storage_1[10][5] ), .B2(n2900), 
        .Z(n3819) );
  aoim22d1 U4652 ( .A1(n2900), .A2(n3053), .B1(\storage_1[10][6] ), .B2(n2900), 
        .Z(n3818) );
  aoim22d1 U4653 ( .A1(n2900), .A2(n3055), .B1(\storage_1[10][7] ), .B2(n2900), 
        .Z(n3817) );
  nd02d0 U4654 ( .A1(n2902), .A2(n2901), .ZN(n2931) );
  nr02d1 U4655 ( .A1(n2903), .A2(n2931), .ZN(n2906) );
  inv0d0 U4656 ( .I(n2906), .ZN(n2905) );
  aoi22d1 U4657 ( .A1(n2906), .A2(n3047), .B1(n2904), .B2(n2905), .ZN(n3816)
         );
  aoim22d1 U4658 ( .A1(n2906), .A2(n3048), .B1(\storage_1[9][1] ), .B2(n2906), 
        .Z(n3815) );
  aoim22d1 U4659 ( .A1(n2906), .A2(n3049), .B1(\storage_1[9][2] ), .B2(n2906), 
        .Z(n3814) );
  aoim22d1 U4660 ( .A1(n2906), .A2(n3050), .B1(\storage_1[9][3] ), .B2(n2906), 
        .Z(n3813) );
  inv0d0 U4661 ( .I(\storage_1[9][4] ), .ZN(n2968) );
  aoi22d1 U4662 ( .A1(n2906), .A2(n3051), .B1(n2968), .B2(n2905), .ZN(n3812)
         );
  aoim22d1 U4663 ( .A1(n2906), .A2(n3052), .B1(\storage_1[9][5] ), .B2(n2906), 
        .Z(n3811) );
  inv0d0 U4664 ( .I(\storage_1[9][6] ), .ZN(n3002) );
  aoi22d1 U4665 ( .A1(n2906), .A2(n3053), .B1(n3002), .B2(n2905), .ZN(n3810)
         );
  aoim22d1 U4666 ( .A1(n2906), .A2(n3055), .B1(\storage_1[9][7] ), .B2(n2906), 
        .Z(n3809) );
  nr02d1 U4667 ( .A1(n2907), .A2(n2931), .ZN(n2908) );
  aoim22d1 U4668 ( .A1(n2908), .A2(n3047), .B1(\storage_1[8][0] ), .B2(n2908), 
        .Z(n3808) );
  aoim22d1 U4669 ( .A1(n2908), .A2(n3048), .B1(\storage_1[8][1] ), .B2(n2908), 
        .Z(n3807) );
  aoim22d1 U4670 ( .A1(n2908), .A2(n3049), .B1(\storage_1[8][2] ), .B2(n2908), 
        .Z(n3806) );
  aoim22d1 U4671 ( .A1(n2908), .A2(n3050), .B1(\storage_1[8][3] ), .B2(n2908), 
        .Z(n3805) );
  aoim22d1 U4672 ( .A1(n2908), .A2(n3051), .B1(\storage_1[8][4] ), .B2(n2908), 
        .Z(n3804) );
  aoim22d1 U4673 ( .A1(n2908), .A2(n3052), .B1(\storage_1[8][5] ), .B2(n2908), 
        .Z(n3803) );
  aoim22d1 U4674 ( .A1(n2908), .A2(n3053), .B1(\storage_1[8][6] ), .B2(n2908), 
        .Z(n3802) );
  aoim22d1 U4675 ( .A1(n2908), .A2(n3055), .B1(\storage_1[8][7] ), .B2(n2908), 
        .Z(n3801) );
  inv0d0 U4676 ( .I(uart_rx_fifo_produce[3]), .ZN(n2914) );
  nd02d0 U4677 ( .A1(n2909), .A2(n2914), .ZN(n2926) );
  nr02d1 U4678 ( .A1(n2916), .A2(n2926), .ZN(n2912) );
  inv0d0 U4679 ( .I(n2912), .ZN(n2911) );
  aoi22d1 U4680 ( .A1(n2912), .A2(n3047), .B1(n2910), .B2(n2911), .ZN(n3800)
         );
  aoim22d1 U4681 ( .A1(n2912), .A2(n3048), .B1(\storage_1[7][1] ), .B2(n2912), 
        .Z(n3799) );
  aoim22d1 U4682 ( .A1(n2912), .A2(n3049), .B1(\storage_1[7][2] ), .B2(n2912), 
        .Z(n3798) );
  aoim22d1 U4683 ( .A1(n2912), .A2(n3050), .B1(\storage_1[7][3] ), .B2(n2912), 
        .Z(n3797) );
  inv0d0 U4684 ( .I(\storage_1[7][4] ), .ZN(n2970) );
  aoi22d1 U4685 ( .A1(n2912), .A2(n3051), .B1(n2970), .B2(n2911), .ZN(n3796)
         );
  aoim22d1 U4686 ( .A1(n2912), .A2(n3052), .B1(\storage_1[7][5] ), .B2(n2912), 
        .Z(n3795) );
  inv0d0 U4687 ( .I(\storage_1[7][6] ), .ZN(n3006) );
  aoi22d1 U4688 ( .A1(n2912), .A2(n3053), .B1(n3006), .B2(n2911), .ZN(n3794)
         );
  aoim22d1 U4689 ( .A1(n2912), .A2(n3055), .B1(\storage_1[7][7] ), .B2(n2912), 
        .Z(n3793) );
  nr02d1 U4690 ( .A1(n2916), .A2(n2930), .ZN(n2917) );
  aoim22d1 U4691 ( .A1(n2917), .A2(n3047), .B1(\storage_1[6][0] ), .B2(n2917), 
        .Z(n3792) );
  aoim22d1 U4692 ( .A1(n2917), .A2(n3048), .B1(\storage_1[6][1] ), .B2(n2917), 
        .Z(n3791) );
  aoim22d1 U4693 ( .A1(n2917), .A2(n3049), .B1(\storage_1[6][2] ), .B2(n2917), 
        .Z(n3790) );
  aoim22d1 U4694 ( .A1(n2917), .A2(n3050), .B1(\storage_1[6][3] ), .B2(n2917), 
        .Z(n3789) );
  aoim22d1 U4695 ( .A1(n2917), .A2(n3051), .B1(\storage_1[6][4] ), .B2(n2917), 
        .Z(n3788) );
  aoim22d1 U4696 ( .A1(n2917), .A2(n3052), .B1(\storage_1[6][5] ), .B2(n2917), 
        .Z(n3787) );
  aoim22d1 U4697 ( .A1(n2917), .A2(n3053), .B1(\storage_1[6][6] ), .B2(n2917), 
        .Z(n3786) );
  aoim22d1 U4698 ( .A1(n2917), .A2(n3055), .B1(\storage_1[6][7] ), .B2(n2917), 
        .Z(n3785) );
  nr02d1 U4699 ( .A1(n2921), .A2(n2926), .ZN(n2920) );
  inv0d0 U4700 ( .I(n2920), .ZN(n2919) );
  aoi22d1 U4701 ( .A1(n2920), .A2(n3047), .B1(n2918), .B2(n2919), .ZN(n3784)
         );
  aoim22d1 U4702 ( .A1(n2920), .A2(n3048), .B1(\storage_1[5][1] ), .B2(n2920), 
        .Z(n3783) );
  aoim22d1 U4703 ( .A1(n2920), .A2(n3049), .B1(\storage_1[5][2] ), .B2(n2920), 
        .Z(n3782) );
  aoim22d1 U4704 ( .A1(n2920), .A2(n3050), .B1(\storage_1[5][3] ), .B2(n2920), 
        .Z(n3781) );
  inv0d0 U4705 ( .I(\storage_1[5][4] ), .ZN(n2967) );
  aoi22d1 U4706 ( .A1(n2920), .A2(n3051), .B1(n2967), .B2(n2919), .ZN(n3780)
         );
  aoim22d1 U4707 ( .A1(n2920), .A2(n3052), .B1(\storage_1[5][5] ), .B2(n2920), 
        .Z(n3779) );
  inv0d0 U4708 ( .I(\storage_1[5][6] ), .ZN(n3000) );
  aoi22d1 U4709 ( .A1(n2920), .A2(n3053), .B1(n3000), .B2(n2919), .ZN(n3778)
         );
  aoim22d1 U4710 ( .A1(n2920), .A2(n3055), .B1(\storage_1[5][7] ), .B2(n2920), 
        .Z(n3777) );
  nr02d1 U4711 ( .A1(n2921), .A2(n2930), .ZN(n2922) );
  aoim22d1 U4712 ( .A1(n2922), .A2(n3047), .B1(\storage_1[4][0] ), .B2(n2922), 
        .Z(n3776) );
  aoim22d1 U4713 ( .A1(n2922), .A2(n3048), .B1(\storage_1[4][1] ), .B2(n2922), 
        .Z(n3775) );
  aoim22d1 U4714 ( .A1(n2922), .A2(n3049), .B1(\storage_1[4][2] ), .B2(n2922), 
        .Z(n3774) );
  aoim22d1 U4715 ( .A1(n2922), .A2(n3050), .B1(\storage_1[4][3] ), .B2(n2922), 
        .Z(n3773) );
  aoim22d1 U4716 ( .A1(n2922), .A2(n3051), .B1(\storage_1[4][4] ), .B2(n2922), 
        .Z(n3772) );
  aoim22d1 U4717 ( .A1(n2922), .A2(n3052), .B1(\storage_1[4][5] ), .B2(n2922), 
        .Z(n3771) );
  aoim22d1 U4718 ( .A1(n2922), .A2(n3053), .B1(\storage_1[4][6] ), .B2(n2922), 
        .Z(n3770) );
  aoim22d1 U4719 ( .A1(n2922), .A2(n3055), .B1(\storage_1[4][7] ), .B2(n2922), 
        .Z(n3769) );
  nr02d1 U4720 ( .A1(n2924), .A2(n2926), .ZN(n2923) );
  aoim22d1 U4721 ( .A1(n2923), .A2(n3047), .B1(\storage_1[3][0] ), .B2(n2923), 
        .Z(n3768) );
  aoim22d1 U4722 ( .A1(n2923), .A2(n3048), .B1(\storage_1[3][1] ), .B2(n2923), 
        .Z(n3767) );
  aoim22d1 U4723 ( .A1(n2923), .A2(n3049), .B1(\storage_1[3][2] ), .B2(n2923), 
        .Z(n3766) );
  aoim22d1 U4724 ( .A1(n2923), .A2(n3050), .B1(\storage_1[3][3] ), .B2(n2923), 
        .Z(n3765) );
  aoim22d1 U4725 ( .A1(n2923), .A2(n3051), .B1(\storage_1[3][4] ), .B2(n2923), 
        .Z(n3764) );
  aoim22d1 U4726 ( .A1(n2923), .A2(n3052), .B1(\storage_1[3][5] ), .B2(n2923), 
        .Z(n3763) );
  aoim22d1 U4727 ( .A1(n2923), .A2(n3053), .B1(\storage_1[3][6] ), .B2(n2923), 
        .Z(n3762) );
  aoim22d1 U4728 ( .A1(n2923), .A2(n3055), .B1(\storage_1[3][7] ), .B2(n2923), 
        .Z(n3761) );
  nr02d1 U4729 ( .A1(n2924), .A2(n2930), .ZN(n2925) );
  aoim22d1 U4730 ( .A1(n2925), .A2(n3047), .B1(\storage_1[2][0] ), .B2(n2925), 
        .Z(n3760) );
  aoim22d1 U4731 ( .A1(n2925), .A2(n3048), .B1(\storage_1[2][1] ), .B2(n2925), 
        .Z(n3759) );
  aoim22d1 U4732 ( .A1(n2925), .A2(n3049), .B1(\storage_1[2][2] ), .B2(n2925), 
        .Z(n3758) );
  aoim22d1 U4733 ( .A1(n2925), .A2(n3050), .B1(\storage_1[2][3] ), .B2(n2925), 
        .Z(n3757) );
  aoim22d1 U4734 ( .A1(n2925), .A2(n3051), .B1(\storage_1[2][4] ), .B2(n2925), 
        .Z(n3756) );
  aoim22d1 U4735 ( .A1(n2925), .A2(n3052), .B1(\storage_1[2][5] ), .B2(n2925), 
        .Z(n3755) );
  aoim22d1 U4736 ( .A1(n2925), .A2(n3053), .B1(\storage_1[2][6] ), .B2(n2925), 
        .Z(n3754) );
  aoim22d1 U4737 ( .A1(n2925), .A2(n3055), .B1(\storage_1[2][7] ), .B2(n2925), 
        .Z(n3753) );
  nr02d1 U4738 ( .A1(n2931), .A2(n2926), .ZN(n2929) );
  inv0d0 U4739 ( .I(n2929), .ZN(n2928) );
  aoi22d1 U4740 ( .A1(n2929), .A2(n3047), .B1(n2927), .B2(n2928), .ZN(n3752)
         );
  aoim22d1 U4741 ( .A1(n2929), .A2(n3048), .B1(\storage_1[1][1] ), .B2(n2929), 
        .Z(n3751) );
  aoim22d1 U4742 ( .A1(n2929), .A2(n3049), .B1(\storage_1[1][2] ), .B2(n2929), 
        .Z(n3750) );
  aoim22d1 U4743 ( .A1(n2929), .A2(n3050), .B1(\storage_1[1][3] ), .B2(n2929), 
        .Z(n3749) );
  inv0d0 U4744 ( .I(\storage_1[1][4] ), .ZN(n2969) );
  aoi22d1 U4745 ( .A1(n2929), .A2(n3051), .B1(n2969), .B2(n2928), .ZN(n3748)
         );
  aoim22d1 U4746 ( .A1(n2929), .A2(n3052), .B1(\storage_1[1][5] ), .B2(n2929), 
        .Z(n3747) );
  inv0d0 U4747 ( .I(\storage_1[1][6] ), .ZN(n2998) );
  aoi22d1 U4748 ( .A1(n2929), .A2(n3053), .B1(n2998), .B2(n2928), .ZN(n3746)
         );
  aoim22d1 U4749 ( .A1(n2929), .A2(n3055), .B1(\storage_1[1][7] ), .B2(n2929), 
        .Z(n3745) );
  nr02d1 U4750 ( .A1(n2931), .A2(n2930), .ZN(n3025) );
  aoim22d1 U4751 ( .A1(n3025), .A2(n3047), .B1(\storage_1[0][0] ), .B2(n3025), 
        .Z(n3744) );
  aoim22d1 U4752 ( .A1(n3025), .A2(n3048), .B1(\storage_1[0][1] ), .B2(n3025), 
        .Z(n3743) );
  aoi22d1 U4753 ( .A1(\storage_1[13][1] ), .A2(n2985), .B1(\storage_1[3][1] ), 
        .B2(n2959), .ZN(n2935) );
  aoi22d1 U4754 ( .A1(\storage_1[15][1] ), .A2(n3033), .B1(\storage_1[9][1] ), 
        .B2(n3013), .ZN(n2934) );
  aoi22d1 U4755 ( .A1(\storage_1[5][1] ), .A2(n3031), .B1(\storage_1[1][1] ), 
        .B2(n2958), .ZN(n2933) );
  aoi22d1 U4756 ( .A1(\storage_1[11][1] ), .A2(n2984), .B1(\storage_1[7][1] ), 
        .B2(n3036), .ZN(n2932) );
  aoi22d1 U4757 ( .A1(\storage_1[4][1] ), .A2(n3031), .B1(\storage_1[2][1] ), 
        .B2(n2959), .ZN(n2939) );
  aoi22d1 U4758 ( .A1(\storage_1[14][1] ), .A2(n3033), .B1(\storage_1[0][1] ), 
        .B2(n2958), .ZN(n2938) );
  aoi22d1 U4759 ( .A1(\storage_1[8][1] ), .A2(n3013), .B1(\storage_1[6][1] ), 
        .B2(n3036), .ZN(n2937) );
  aoi22d1 U4760 ( .A1(\storage_1[12][1] ), .A2(n2985), .B1(\storage_1[10][1] ), 
        .B2(n3035), .ZN(n2936) );
  aoi22d1 U4761 ( .A1(uart_rx_fifo_rdport_adr[0]), .A2(n2941), .B1(n2940), 
        .B2(n3042), .ZN(n2942) );
  aoim22d1 U4762 ( .A1(n3046), .A2(n2942), .B1(
        uart_rx_fifo_fifo_out_payload_data[1]), .B2(n3046), .Z(n3742) );
  aoim22d1 U4763 ( .A1(n3025), .A2(n3049), .B1(\storage_1[0][2] ), .B2(n3025), 
        .Z(n3741) );
  aoi22d1 U4764 ( .A1(\storage_1[7][2] ), .A2(n3036), .B1(\storage_1[1][2] ), 
        .B2(n2958), .ZN(n2946) );
  aoi22d1 U4765 ( .A1(\storage_1[11][2] ), .A2(n2984), .B1(\storage_1[3][2] ), 
        .B2(n2959), .ZN(n2945) );
  aoi22d1 U4766 ( .A1(\storage_1[15][2] ), .A2(n3033), .B1(\storage_1[13][2] ), 
        .B2(n3037), .ZN(n2944) );
  aoi22d1 U4767 ( .A1(\storage_1[9][2] ), .A2(n3013), .B1(\storage_1[5][2] ), 
        .B2(n3012), .ZN(n2943) );
  aoi22d1 U4768 ( .A1(\storage_1[10][2] ), .A2(n3035), .B1(\storage_1[0][2] ), 
        .B2(n2958), .ZN(n2950) );
  aoi22d1 U4769 ( .A1(\storage_1[12][2] ), .A2(n2985), .B1(\storage_1[8][2] ), 
        .B2(n3034), .ZN(n2949) );
  aoi22d1 U4770 ( .A1(\storage_1[6][2] ), .A2(n3036), .B1(\storage_1[4][2] ), 
        .B2(n3012), .ZN(n2948) );
  aoi22d1 U4771 ( .A1(\storage_1[14][2] ), .A2(n3033), .B1(\storage_1[2][2] ), 
        .B2(n2959), .ZN(n2947) );
  aoi22d1 U4772 ( .A1(uart_rx_fifo_rdport_adr[0]), .A2(n2952), .B1(n2951), 
        .B2(n3042), .ZN(n2953) );
  aoim22d1 U4773 ( .A1(n3046), .A2(n2953), .B1(
        uart_rx_fifo_fifo_out_payload_data[2]), .B2(n3046), .Z(n3740) );
  aoim22d1 U4774 ( .A1(n3025), .A2(n3050), .B1(\storage_1[0][3] ), .B2(n3025), 
        .Z(n3739) );
  aoi22d1 U4775 ( .A1(\storage_1[11][3] ), .A2(n2984), .B1(\storage_1[7][3] ), 
        .B2(n3036), .ZN(n2957) );
  aoi22d1 U4776 ( .A1(\storage_1[15][3] ), .A2(n3033), .B1(\storage_1[3][3] ), 
        .B2(n2959), .ZN(n2956) );
  aoi22d1 U4777 ( .A1(\storage_1[13][3] ), .A2(n2985), .B1(\storage_1[9][3] ), 
        .B2(n3034), .ZN(n2955) );
  aoi22d1 U4778 ( .A1(\storage_1[5][3] ), .A2(n3031), .B1(\storage_1[1][3] ), 
        .B2(n2958), .ZN(n2954) );
  aoi22d1 U4779 ( .A1(\storage_1[6][3] ), .A2(n3036), .B1(\storage_1[4][3] ), 
        .B2(n3012), .ZN(n2963) );
  aoi22d1 U4780 ( .A1(\storage_1[2][3] ), .A2(n2959), .B1(\storage_1[0][3] ), 
        .B2(n2958), .ZN(n2962) );
  aoi22d1 U4781 ( .A1(\storage_1[14][3] ), .A2(n3033), .B1(\storage_1[12][3] ), 
        .B2(n3037), .ZN(n2961) );
  aoi22d1 U4782 ( .A1(\storage_1[10][3] ), .A2(n2984), .B1(\storage_1[8][3] ), 
        .B2(n3034), .ZN(n2960) );
  aoi22d1 U4783 ( .A1(uart_rx_fifo_rdport_adr[0]), .A2(n2965), .B1(n2964), 
        .B2(n3042), .ZN(n2966) );
  aoim22d1 U4784 ( .A1(n3046), .A2(n2966), .B1(
        uart_rx_fifo_fifo_out_payload_data[3]), .B2(n3046), .Z(n3738) );
  aoim22d1 U4785 ( .A1(n3025), .A2(n3051), .B1(\storage_1[0][4] ), .B2(n3025), 
        .Z(n3737) );
  aoi22d1 U4786 ( .A1(\storage_1[11][4] ), .A2(n2984), .B1(\storage_1[3][4] ), 
        .B2(n3032), .ZN(n2983) );
  oai22d1 U4787 ( .A1(n2968), .A2(n3001), .B1(n2967), .B2(n2999), .ZN(n2975)
         );
  oai22d1 U4788 ( .A1(n2970), .A2(n3005), .B1(n2969), .B2(n2997), .ZN(n2974)
         );
  oai22d1 U4789 ( .A1(n2972), .A2(n3003), .B1(n2971), .B2(n3007), .ZN(n2973)
         );
  aoi22d1 U4790 ( .A1(\storage_1[12][4] ), .A2(n2985), .B1(\storage_1[10][4] ), 
        .B2(n3035), .ZN(n2979) );
  aoi22d1 U4791 ( .A1(\storage_1[14][4] ), .A2(n3033), .B1(\storage_1[8][4] ), 
        .B2(n3034), .ZN(n2978) );
  aoi22d1 U4792 ( .A1(\storage_1[6][4] ), .A2(n3036), .B1(\storage_1[0][4] ), 
        .B2(n3030), .ZN(n2977) );
  aoi22d1 U4793 ( .A1(\storage_1[4][4] ), .A2(n3031), .B1(\storage_1[2][4] ), 
        .B2(n3032), .ZN(n2976) );
  aoi22d1 U4794 ( .A1(uart_rx_fifo_fifo_out_payload_data[4]), .A2(n3020), .B1(
        n3019), .B2(n2980), .ZN(n2981) );
  aon211d1 U4795 ( .C1(n2983), .C2(n2982), .B(n3022), .A(n2981), .ZN(n3736) );
  aoim22d1 U4796 ( .A1(n3025), .A2(n3052), .B1(\storage_1[0][5] ), .B2(n3025), 
        .Z(n3735) );
  aoi22d1 U4797 ( .A1(\storage_1[9][5] ), .A2(n3013), .B1(\storage_1[3][5] ), 
        .B2(n3032), .ZN(n2989) );
  aoi22d1 U4798 ( .A1(\storage_1[11][5] ), .A2(n2984), .B1(\storage_1[5][5] ), 
        .B2(n3012), .ZN(n2988) );
  aoi22d1 U4799 ( .A1(\storage_1[13][5] ), .A2(n2985), .B1(\storage_1[7][5] ), 
        .B2(n3036), .ZN(n2987) );
  aoi22d1 U4800 ( .A1(\storage_1[15][5] ), .A2(n3033), .B1(\storage_1[1][5] ), 
        .B2(n3030), .ZN(n2986) );
  aoi22d1 U4801 ( .A1(\storage_1[8][5] ), .A2(n3013), .B1(\storage_1[2][5] ), 
        .B2(n3032), .ZN(n2993) );
  aoi22d1 U4802 ( .A1(\storage_1[14][5] ), .A2(n3033), .B1(\storage_1[12][5] ), 
        .B2(n3037), .ZN(n2992) );
  aoi22d1 U4803 ( .A1(\storage_1[6][5] ), .A2(n3036), .B1(\storage_1[4][5] ), 
        .B2(n3012), .ZN(n2991) );
  aoi22d1 U4804 ( .A1(\storage_1[10][5] ), .A2(n3035), .B1(\storage_1[0][5] ), 
        .B2(n3030), .ZN(n2990) );
  aoi22d1 U4805 ( .A1(uart_rx_fifo_rdport_adr[0]), .A2(n2995), .B1(n2994), 
        .B2(n3042), .ZN(n2996) );
  aoim22d1 U4806 ( .A1(n3046), .A2(n2996), .B1(
        uart_rx_fifo_fifo_out_payload_data[5]), .B2(n3046), .Z(n3734) );
  aoim22d1 U4807 ( .A1(n3025), .A2(n3053), .B1(\storage_1[0][6] ), .B2(n3025), 
        .Z(n3733) );
  aoi22d1 U4808 ( .A1(\storage_1[11][6] ), .A2(n3035), .B1(\storage_1[3][6] ), 
        .B2(n3032), .ZN(n3024) );
  oai22d1 U4809 ( .A1(n3000), .A2(n2999), .B1(n2998), .B2(n2997), .ZN(n3011)
         );
  oai22d1 U4810 ( .A1(n3004), .A2(n3003), .B1(n3002), .B2(n3001), .ZN(n3010)
         );
  oai22d1 U4811 ( .A1(n3008), .A2(n3007), .B1(n3006), .B2(n3005), .ZN(n3009)
         );
  aoi22d1 U4812 ( .A1(\storage_1[14][6] ), .A2(n3033), .B1(\storage_1[6][6] ), 
        .B2(n3036), .ZN(n3017) );
  aoi22d1 U4813 ( .A1(\storage_1[10][6] ), .A2(n3035), .B1(\storage_1[2][6] ), 
        .B2(n3032), .ZN(n3016) );
  aoi22d1 U4814 ( .A1(\storage_1[12][6] ), .A2(n3037), .B1(\storage_1[4][6] ), 
        .B2(n3012), .ZN(n3015) );
  aoi22d1 U4815 ( .A1(\storage_1[8][6] ), .A2(n3013), .B1(\storage_1[0][6] ), 
        .B2(n3030), .ZN(n3014) );
  aoi22d1 U4816 ( .A1(uart_rx_fifo_fifo_out_payload_data[6]), .A2(n3020), .B1(
        n3019), .B2(n3018), .ZN(n3021) );
  aon211d1 U4817 ( .C1(n3024), .C2(n3023), .B(n3022), .A(n3021), .ZN(n3732) );
  aoim22d1 U4818 ( .A1(n3025), .A2(n3055), .B1(\storage_1[0][7] ), .B2(n3025), 
        .Z(n3731) );
  aoi22d1 U4819 ( .A1(\storage_1[13][7] ), .A2(n3037), .B1(\storage_1[9][7] ), 
        .B2(n3034), .ZN(n3029) );
  aoi22d1 U4820 ( .A1(\storage_1[15][7] ), .A2(n3033), .B1(\storage_1[1][7] ), 
        .B2(n3030), .ZN(n3028) );
  aoi22d1 U4821 ( .A1(\storage_1[5][7] ), .A2(n3031), .B1(\storage_1[3][7] ), 
        .B2(n3032), .ZN(n3027) );
  aoi22d1 U4822 ( .A1(\storage_1[11][7] ), .A2(n3035), .B1(\storage_1[7][7] ), 
        .B2(n3036), .ZN(n3026) );
  aoi22d1 U4823 ( .A1(\storage_1[4][7] ), .A2(n3031), .B1(\storage_1[0][7] ), 
        .B2(n3030), .ZN(n3041) );
  aoi22d1 U4824 ( .A1(\storage_1[14][7] ), .A2(n3033), .B1(\storage_1[2][7] ), 
        .B2(n3032), .ZN(n3040) );
  aoi22d1 U4825 ( .A1(\storage_1[10][7] ), .A2(n3035), .B1(\storage_1[8][7] ), 
        .B2(n3034), .ZN(n3039) );
  aoi22d1 U4826 ( .A1(\storage_1[12][7] ), .A2(n3037), .B1(\storage_1[6][7] ), 
        .B2(n3036), .ZN(n3038) );
  aoi22d1 U4827 ( .A1(uart_rx_fifo_rdport_adr[0]), .A2(n3044), .B1(n3043), 
        .B2(n3042), .ZN(n3045) );
  aoim22d1 U4828 ( .A1(n3046), .A2(n3045), .B1(
        uart_rx_fifo_fifo_out_payload_data[7]), .B2(n3046), .Z(n3730) );
  aoi22d1 U4829 ( .A1(n3057), .A2(n3048), .B1(n3047), .B2(n3054), .ZN(n3729)
         );
  aoi22d1 U4830 ( .A1(n3057), .A2(n3049), .B1(n3048), .B2(n3054), .ZN(n3728)
         );
  aoi22d1 U4831 ( .A1(n3057), .A2(n3050), .B1(n3049), .B2(n3054), .ZN(n3727)
         );
  aoi22d1 U4832 ( .A1(n3057), .A2(n3051), .B1(n3050), .B2(n3054), .ZN(n3726)
         );
  aoi22d1 U4833 ( .A1(n3057), .A2(n3053), .B1(n3052), .B2(n3054), .ZN(n3724)
         );
  aoi22d1 U4834 ( .A1(n3057), .A2(n3055), .B1(n3053), .B2(n3054), .ZN(n3723)
         );
  aoi22d1 U4835 ( .A1(n3057), .A2(n3056), .B1(n3055), .B2(n3054), .ZN(n3722)
         );
  nr04d0 U4836 ( .A1(n4811), .A2(n3060), .A3(n3059), .A4(n3058), .ZN(n3062) );
  oai21d1 U4837 ( .B1(mprj_wb_iena), .B2(n3062), .A(n5319), .ZN(n3061) );
  aoi21d1 U4838 ( .B1(n3062), .B2(n4808), .A(n3061), .ZN(n3721) );
  nd02d1 U4839 ( .A1(n4580), .A2(n3063), .ZN(n3081) );
  nd02d1 U4840 ( .A1(n5955), .A2(n3081), .ZN(n3080) );
  inv0d0 U4841 ( .I(n3080), .ZN(n3070) );
  oaim22d1 U4842 ( .A1(n5290), .A2(n3081), .B1(n3070), .B2(
        spi_master_clk_divider0[0]), .ZN(n3720) );
  oai22d1 U4843 ( .A1(n5294), .A2(n3081), .B1(n3064), .B2(n3080), .ZN(n3719)
         );
  inv0d0 U4844 ( .I(n3081), .ZN(n3069) );
  aoi22d1 U4845 ( .A1(n3070), .A2(n3065), .B1(n3069), .B2(n5245), .ZN(n3718)
         );
  oai22d1 U4846 ( .A1(n5006), .A2(n3081), .B1(n3066), .B2(n3080), .ZN(n3717)
         );
  oai22d1 U4847 ( .A1(n5008), .A2(n3081), .B1(n3067), .B2(n3080), .ZN(n3716)
         );
  aoi22d1 U4848 ( .A1(n3070), .A2(n3068), .B1(n3069), .B2(n5010), .ZN(n3715)
         );
  aoim22d1 U4849 ( .A1(n3069), .A2(n5012), .B1(n3080), .B2(
        spi_master_clk_divider0[6]), .Z(n3714) );
  oaim22d1 U4850 ( .A1(n3071), .A2(n3081), .B1(spi_master_clk_divider0[7]), 
        .B2(n3070), .ZN(n3713) );
  oai22d1 U4851 ( .A1(n4783), .A2(n3081), .B1(n3080), .B2(n3072), .ZN(n3712)
         );
  oai22d1 U4852 ( .A1(n4593), .A2(n3081), .B1(n3080), .B2(n3073), .ZN(n3711)
         );
  oai22d1 U4853 ( .A1(n4595), .A2(n3081), .B1(n3080), .B2(n3074), .ZN(n3710)
         );
  oai22d1 U4854 ( .A1(n4787), .A2(n3081), .B1(n3080), .B2(n3075), .ZN(n3709)
         );
  oai22d1 U4855 ( .A1(n4598), .A2(n3081), .B1(n3080), .B2(n3076), .ZN(n3708)
         );
  oai22d1 U4856 ( .A1(n4790), .A2(n3081), .B1(n3080), .B2(n3077), .ZN(n3707)
         );
  oai22d1 U4857 ( .A1(n4601), .A2(n3081), .B1(n3080), .B2(n3078), .ZN(n3706)
         );
  oai22d1 U4858 ( .A1(n4793), .A2(n3081), .B1(n3080), .B2(n3079), .ZN(n3705)
         );
  nr02d0 U4859 ( .A1(n5100), .A2(n4679), .ZN(n4623) );
  inv0d0 U4860 ( .I(n4623), .ZN(n3084) );
  inv0d0 U4861 ( .I(spi_master_miso_data[0]), .ZN(n4645) );
  inv0d0 U4862 ( .I(spi_master_loopback), .ZN(n3082) );
  aoi22d1 U4863 ( .A1(spi_master_loopback), .A2(spi_mosi), .B1(spi_miso), .B2(
        n3082), .ZN(n3083) );
  oai22d1 U4864 ( .A1(n3084), .A2(n4645), .B1(n4682), .B2(n3083), .ZN(n3704)
         );
  inv0d0 U4865 ( .I(spi_master_miso_data[1]), .ZN(n4647) );
  oai22d1 U4866 ( .A1(n3084), .A2(n4647), .B1(n4682), .B2(n4645), .ZN(n3703)
         );
  inv0d0 U4867 ( .I(spi_master_miso_data[2]), .ZN(n4649) );
  oai22d1 U4868 ( .A1(n3084), .A2(n4649), .B1(n4682), .B2(n4647), .ZN(n3702)
         );
  inv0d0 U4869 ( .I(spi_master_miso_data[3]), .ZN(n4651) );
  oai22d1 U4870 ( .A1(n3084), .A2(n4651), .B1(n4682), .B2(n4649), .ZN(n3701)
         );
  inv0d0 U4871 ( .I(spi_master_miso_data[4]), .ZN(n4653) );
  oai22d1 U4872 ( .A1(n3084), .A2(n4653), .B1(n4682), .B2(n4651), .ZN(n3700)
         );
  inv0d0 U4873 ( .I(spi_master_miso_data[5]), .ZN(n4655) );
  oai22d1 U4874 ( .A1(n3084), .A2(n4655), .B1(n4682), .B2(n4653), .ZN(n3699)
         );
  inv0d0 U4875 ( .I(spi_master_miso_data[6]), .ZN(n4657) );
  oai22d1 U4876 ( .A1(n3084), .A2(n4657), .B1(n4682), .B2(n4655), .ZN(n3698)
         );
  inv0d0 U4877 ( .I(spi_master_miso_data[7]), .ZN(n4659) );
  oai22d1 U4878 ( .A1(n3084), .A2(n4659), .B1(n4682), .B2(n4657), .ZN(n3697)
         );
  inv0d0 U4879 ( .I(spi_master_mosi_sel[0]), .ZN(n4548) );
  nd03d0 U4880 ( .A1(csrbank9_control0_w[0]), .A2(n3085), .A3(
        spi_master_control_re), .ZN(n4551) );
  nr02d0 U4881 ( .A1(n3089), .A2(n5100), .ZN(n4568) );
  nd02d0 U4882 ( .A1(n4568), .A2(n4548), .ZN(n3086) );
  oai211d1 U4883 ( .C1(n3087), .C2(n4548), .A(n4566), .B(n3086), .ZN(n3696) );
  oai21d1 U4884 ( .B1(spi_master_mosi_sel[0]), .B2(n3089), .A(n5319), .ZN(
        n4550) );
  inv0d0 U4885 ( .I(spi_master_mosi_sel[1]), .ZN(n3119) );
  aoi31d1 U4886 ( .B1(n4568), .B2(n3119), .B3(n4548), .A(n4620), .ZN(n3118) );
  oai21d1 U4887 ( .B1(n4550), .B2(n3119), .A(n3118), .ZN(n3695) );
  inv0d0 U4888 ( .I(spi_master_mosi_sel[2]), .ZN(n4663) );
  nr02d0 U4889 ( .A1(spi_master_mosi_sel[2]), .A2(spi_master_mosi_sel[1]), 
        .ZN(n4669) );
  nr02d0 U4890 ( .A1(n4663), .A2(n3119), .ZN(n4664) );
  aon211d1 U4891 ( .C1(n4669), .C2(n4548), .B(n4664), .A(n4568), .ZN(n4549) );
  oai211d1 U4892 ( .C1(n4550), .C2(n4663), .A(n4549), .B(n4566), .ZN(n3694) );
  inv0d0 U4893 ( .I(spi_master_mosi_data[0]), .ZN(n4552) );
  nd02d0 U4894 ( .A1(n5955), .A2(n4551), .ZN(n4564) );
  oai22d1 U4895 ( .A1(n4553), .A2(n4566), .B1(n4552), .B2(n4564), .ZN(n3693)
         );
  inv0d0 U4896 ( .I(spi_master_mosi_data[1]), .ZN(n4554) );
  oai22d1 U4897 ( .A1(n4555), .A2(n4566), .B1(n4554), .B2(n4564), .ZN(n3692)
         );
  inv0d0 U4898 ( .I(spi_master_mosi_data[2]), .ZN(n4667) );
  oai22d1 U4899 ( .A1(n4556), .A2(n4566), .B1(n4667), .B2(n4564), .ZN(n3691)
         );
  inv0d0 U4900 ( .I(spi_master_mosi_data[3]), .ZN(n4666) );
  oai22d1 U4901 ( .A1(n4557), .A2(n4566), .B1(n4666), .B2(n4564), .ZN(n3690)
         );
  inv0d0 U4902 ( .I(spi_master_mosi_data[4]), .ZN(n4558) );
  oai22d1 U4903 ( .A1(n4559), .A2(n4566), .B1(n4558), .B2(n4564), .ZN(n3689)
         );
  inv0d0 U4904 ( .I(spi_master_mosi_data[5]), .ZN(n4560) );
  oai22d1 U4905 ( .A1(n4561), .A2(n4566), .B1(n4560), .B2(n4564), .ZN(n3688)
         );
  inv0d0 U4906 ( .I(spi_master_mosi_data[6]), .ZN(n4562) );
  oai22d1 U4907 ( .A1(n4563), .A2(n4566), .B1(n4562), .B2(n4564), .ZN(n3687)
         );
  inv0d0 U4908 ( .I(spi_master_mosi_data[7]), .ZN(n4565) );
  oai22d1 U4909 ( .A1(n4567), .A2(n4566), .B1(n4565), .B2(n4564), .ZN(n3686)
         );
  nd02d0 U4910 ( .A1(spimaster_state[1]), .A2(n4625), .ZN(n4681) );
  nd12d0 U4911 ( .A1(n4681), .A2(n4568), .ZN(n4570) );
  inv0d0 U4912 ( .I(spi_master_count[0]), .ZN(n4571) );
  inv0d0 U4913 ( .I(n4570), .ZN(n4572) );
  aoi211d1 U4914 ( .C1(spimaster_state[0]), .C2(n4627), .A(sys_rst), .B(n4572), 
        .ZN(n4569) );
  aoim22d1 U4915 ( .A1(n4570), .A2(n4571), .B1(n4571), .B2(n4569), .Z(n3685)
         );
  inv0d0 U4916 ( .I(spi_master_count[1]), .ZN(n4610) );
  oan211d1 U4917 ( .C1(n4610), .C2(n4571), .B(n4572), .A(n4569), .ZN(n4574) );
  oan211d1 U4918 ( .C1(n4571), .C2(n4570), .B(n4610), .A(n4574), .ZN(n3684) );
  inv0d0 U4919 ( .I(spi_master_count[2]), .ZN(n4607) );
  oai21d1 U4920 ( .B1(n4574), .B2(n4607), .A(n4573), .ZN(n3683) );
  oai21d1 U4921 ( .B1(spi_master_loopback), .B2(n4578), .A(n5955), .ZN(n4577)
         );
  aoi21d1 U4922 ( .B1(n4578), .B2(n5290), .A(n4577), .ZN(n3682) );
  oai22d1 U4923 ( .A1(n4604), .A2(csrbank9_cs0_w[0]), .B1(n4581), .B2(n4582), 
        .ZN(n4583) );
  inv0d0 U4924 ( .I(n4583), .ZN(n3681) );
  inv0d0 U4925 ( .I(csrbank9_cs0_w[1]), .ZN(n4584) );
  oai22d1 U4926 ( .A1(n5294), .A2(n4581), .B1(n4584), .B2(n4604), .ZN(n3680)
         );
  inv0d0 U4927 ( .I(csrbank9_cs0_w[2]), .ZN(n4585) );
  oai22d1 U4928 ( .A1(n5245), .A2(n4581), .B1(n4585), .B2(n4604), .ZN(n3679)
         );
  inv0d0 U4929 ( .I(csrbank9_cs0_w[3]), .ZN(n4586) );
  oai22d1 U4930 ( .A1(n5006), .A2(n4581), .B1(n4586), .B2(n4604), .ZN(n3678)
         );
  inv0d0 U4931 ( .I(csrbank9_cs0_w[4]), .ZN(n4587) );
  oai22d1 U4932 ( .A1(n5008), .A2(n4581), .B1(n4587), .B2(n4604), .ZN(n3677)
         );
  inv0d0 U4933 ( .I(csrbank9_cs0_w[5]), .ZN(n4588) );
  oai22d1 U4934 ( .A1(n5010), .A2(n4581), .B1(n4588), .B2(n4604), .ZN(n3676)
         );
  inv0d0 U4935 ( .I(csrbank9_cs0_w[6]), .ZN(n4589) );
  oai22d1 U4936 ( .A1(n5012), .A2(n4581), .B1(n4589), .B2(n4604), .ZN(n3675)
         );
  inv0d0 U4937 ( .I(csrbank9_cs0_w[7]), .ZN(n4590) );
  oai22d1 U4938 ( .A1(n5251), .A2(n4581), .B1(n4590), .B2(n4604), .ZN(n3674)
         );
  oai22d1 U4939 ( .A1(n5015), .A2(n4581), .B1(n4604), .B2(n4591), .ZN(n3673)
         );
  oai22d1 U4940 ( .A1(n4593), .A2(n4581), .B1(n4604), .B2(n4592), .ZN(n3672)
         );
  oai22d1 U4941 ( .A1(n4595), .A2(n4581), .B1(n4604), .B2(n4594), .ZN(n3671)
         );
  oai22d1 U4942 ( .A1(n4787), .A2(n4581), .B1(n4604), .B2(n4596), .ZN(n3670)
         );
  oai22d1 U4943 ( .A1(n4598), .A2(n4581), .B1(n4604), .B2(n4597), .ZN(n3669)
         );
  oai22d1 U4944 ( .A1(n5024), .A2(n4581), .B1(n4604), .B2(n4599), .ZN(n3668)
         );
  oai22d1 U4945 ( .A1(n4601), .A2(n4581), .B1(n4604), .B2(n4600), .ZN(n3667)
         );
  oai22d1 U4946 ( .A1(n5028), .A2(n4581), .B1(n4604), .B2(n4602), .ZN(n3666)
         );
  oai22d1 U4947 ( .A1(n2003), .A2(n4581), .B1(n4604), .B2(n4603), .ZN(n3665)
         );
  inv0d1 U4948 ( .I(N5618), .ZN(n4644) );
  nd02d1 U4949 ( .A1(n5955), .A2(n4644), .ZN(n4643) );
  inv0d0 U4950 ( .I(csrbank9_control0_w[0]), .ZN(n4605) );
  oai22d1 U4951 ( .A1(n4808), .A2(n4644), .B1(n4643), .B2(n4605), .ZN(n3664)
         );
  nd02d0 U4952 ( .A1(spi_master_count[1]), .A2(n4636), .ZN(n4612) );
  nd02d0 U4953 ( .A1(spi_master_count[2]), .A2(n4638), .ZN(n4606) );
  oan211d1 U4954 ( .C1(spi_master_count[2]), .C2(n4612), .B(n4606), .A(
        spi_master_length0[2]), .ZN(n4619) );
  oan211d1 U4955 ( .C1(spi_master_count[1]), .C2(n4636), .B(
        spi_master_length0[0]), .A(spi_master_count[0]), .ZN(n4618) );
  inv0d0 U4956 ( .I(n4612), .ZN(n4608) );
  nd02d0 U4957 ( .A1(n4635), .A2(n4636), .ZN(n4609) );
  aoi221d1 U4958 ( .B1(spi_master_count[2]), .B2(n4608), .C1(n4607), .C2(n4609), .A(spi_master_length0[3]), .ZN(n4615) );
  aoi211d1 U4959 ( .C1(spi_master_length0[3]), .C2(n4609), .A(
        spi_master_length0[4]), .B(n4681), .ZN(n4614) );
  nd02d0 U4960 ( .A1(spi_master_length0[1]), .A2(n4610), .ZN(n4611) );
  aon211d1 U4961 ( .C1(n4612), .C2(n4611), .B(spi_master_length0[0]), .A(
        spi_master_count[0]), .ZN(n4613) );
  oai211d1 U4962 ( .C1(n4637), .C2(n4615), .A(n4614), .B(n4613), .ZN(n4616) );
  nr04d0 U4963 ( .A1(n4619), .A2(n4618), .A3(n4617), .A4(n4616), .ZN(n4621) );
  aoi211d1 U4964 ( .C1(n4623), .C2(n4622), .A(n4621), .B(n4620), .ZN(n4624) );
  aoi31d1 U4965 ( .B1(n4678), .B2(spimaster_state[1]), .B3(n4625), .A(n4624), 
        .ZN(n4626) );
  aor31d1 U4966 ( .B1(n4678), .B2(spimaster_state[0]), .B3(n4627), .A(n4626), 
        .Z(n3662) );
  inv0d0 U4967 ( .I(csrbank9_control0_w[1]), .ZN(n4628) );
  oai22d1 U4968 ( .A1(n5294), .A2(n4644), .B1(n4628), .B2(n4643), .ZN(n3661)
         );
  inv0d0 U4969 ( .I(csrbank9_control0_w[2]), .ZN(n4629) );
  oai22d1 U4970 ( .A1(n5245), .A2(n4644), .B1(n4629), .B2(n4643), .ZN(n3660)
         );
  inv0d0 U4971 ( .I(csrbank9_control0_w[3]), .ZN(n4630) );
  oai22d1 U4972 ( .A1(n5006), .A2(n4644), .B1(n4630), .B2(n4643), .ZN(n3659)
         );
  inv0d0 U4973 ( .I(csrbank9_control0_w[4]), .ZN(n4631) );
  oai22d1 U4974 ( .A1(n5008), .A2(n4644), .B1(n4631), .B2(n4643), .ZN(n3658)
         );
  inv0d0 U4975 ( .I(csrbank9_control0_w[5]), .ZN(n4632) );
  oai22d1 U4976 ( .A1(n5010), .A2(n4644), .B1(n4632), .B2(n4643), .ZN(n3657)
         );
  inv0d0 U4977 ( .I(csrbank9_control0_w[6]), .ZN(n4633) );
  oai22d1 U4978 ( .A1(n5012), .A2(n4644), .B1(n4633), .B2(n4643), .ZN(n3656)
         );
  inv0d0 U4979 ( .I(csrbank9_control0_w[7]), .ZN(n4634) );
  oai22d1 U4980 ( .A1(n5251), .A2(n4644), .B1(n4634), .B2(n4643), .ZN(n3655)
         );
  oai22d1 U4981 ( .A1(n4783), .A2(n4644), .B1(n4643), .B2(n4635), .ZN(n3654)
         );
  oai22d1 U4982 ( .A1(n4593), .A2(n4644), .B1(n4643), .B2(n4636), .ZN(n3653)
         );
  oai22d1 U4983 ( .A1(n4595), .A2(n4644), .B1(n4643), .B2(n4637), .ZN(n3652)
         );
  oai22d1 U4984 ( .A1(n5254), .A2(n4644), .B1(n4643), .B2(n4638), .ZN(n3651)
         );
  oai22d1 U4985 ( .A1(n4598), .A2(n4644), .B1(n4643), .B2(n4639), .ZN(n3650)
         );
  oai22d1 U4986 ( .A1(n4790), .A2(n4644), .B1(n4643), .B2(n4640), .ZN(n3649)
         );
  oai22d1 U4987 ( .A1(n4601), .A2(n4644), .B1(n4643), .B2(n4641), .ZN(n3648)
         );
  oai22d1 U4988 ( .A1(n4793), .A2(n4644), .B1(n4643), .B2(n4642), .ZN(n3647)
         );
  inv0d0 U4989 ( .I(spi_master_miso_status[0]), .ZN(n4646) );
  oai22d1 U4990 ( .A1(n4646), .A2(n4661), .B1(n4660), .B2(n4645), .ZN(n3646)
         );
  inv0d0 U4991 ( .I(spi_master_miso_status[1]), .ZN(n4648) );
  oai22d1 U4992 ( .A1(n4648), .A2(n4661), .B1(n4660), .B2(n4647), .ZN(n3645)
         );
  inv0d0 U4993 ( .I(spi_master_miso_status[2]), .ZN(n4650) );
  oai22d1 U4994 ( .A1(n4650), .A2(n4661), .B1(n4660), .B2(n4649), .ZN(n3644)
         );
  inv0d0 U4995 ( .I(spi_master_miso_status[3]), .ZN(n4652) );
  oai22d1 U4996 ( .A1(n4652), .A2(n4661), .B1(n4660), .B2(n4651), .ZN(n3643)
         );
  inv0d0 U4997 ( .I(spi_master_miso_status[4]), .ZN(n4654) );
  oai22d1 U4998 ( .A1(n4654), .A2(n4661), .B1(n4660), .B2(n4653), .ZN(n3642)
         );
  inv0d0 U4999 ( .I(spi_master_miso_status[5]), .ZN(n4656) );
  oai22d1 U5000 ( .A1(n4656), .A2(n4661), .B1(n4660), .B2(n4655), .ZN(n3641)
         );
  inv0d0 U5001 ( .I(spi_master_miso_status[6]), .ZN(n4658) );
  oai22d1 U5002 ( .A1(n4658), .A2(n4661), .B1(n4660), .B2(n4657), .ZN(n3640)
         );
  inv0d0 U5003 ( .I(spi_master_miso_status[7]), .ZN(n4662) );
  oai22d1 U5004 ( .A1(n4662), .A2(n4661), .B1(n4660), .B2(n4659), .ZN(n3639)
         );
  nr02d0 U5005 ( .A1(spi_master_mosi_sel[1]), .A2(n4663), .ZN(n4674) );
  nd02d0 U5006 ( .A1(spi_master_mosi_sel[1]), .A2(n4663), .ZN(n4668) );
  aoi22d1 U5007 ( .A1(n4669), .A2(spi_master_mosi_data[1]), .B1(n4664), .B2(
        spi_master_mosi_data[7]), .ZN(n4665) );
  oai211d1 U5008 ( .C1(n4668), .C2(n4666), .A(spi_master_mosi_sel[0]), .B(
        n4665), .ZN(n4673) );
  aoi31d1 U5009 ( .B1(spi_master_mosi_sel[1]), .B2(spi_master_mosi_sel[2]), 
        .B3(spi_master_mosi_data[6]), .A(spi_master_mosi_sel[0]), .ZN(n4671)
         );
  aoim22d1 U5010 ( .A1(n4669), .A2(spi_master_mosi_data[0]), .B1(n4668), .B2(
        n4667), .Z(n4670) );
  oaim211d1 U5011 ( .C1(n4674), .C2(spi_master_mosi_data[4]), .A(n4671), .B(
        n4670), .ZN(n4672) );
  aon211d1 U5012 ( .C1(spi_master_mosi_data[5]), .C2(n4674), .B(n4673), .A(
        n4672), .ZN(n4676) );
  oai21d1 U5013 ( .B1(spi_mosi), .B2(n4677), .A(n5955), .ZN(n4675) );
  aoi21d1 U5014 ( .B1(n4677), .B2(n4676), .A(n4675), .ZN(n3638) );
  nd13d1 U5015 ( .A1(n4679), .A2(n4678), .A3(spi_clk), .ZN(n4680) );
  oai21d1 U5016 ( .B1(n4682), .B2(n4681), .A(n4680), .ZN(n3637) );
  oai211d1 U5017 ( .C1(n4683), .C2(n4723), .A(
        \mgmtsoc_master_status_status[1] ), .B(n4881), .ZN(n4721) );
  buffd1 U5018 ( .I(n4721), .Z(n4717) );
  oai31d1 U5019 ( .B1(n5111), .B2(n4685), .B3(n4684), .A(n4717), .ZN(n3636) );
  inv0d0 U5020 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[0]), .ZN(
        n5739) );
  nd02d1 U5021 ( .A1(n4686), .A2(n5956), .ZN(n4722) );
  buffd1 U5022 ( .I(n4722), .Z(n4718) );
  oai22d1 U5023 ( .A1(n5739), .A2(n4718), .B1(n4717), .B2(n4687), .ZN(n3635)
         );
  inv0d0 U5024 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[1]), .ZN(
        n5740) );
  inv0d0 U5025 ( .I(mgmtsoc_master_rxtx_w[1]), .ZN(n4688) );
  oai22d1 U5026 ( .A1(n4718), .A2(n5740), .B1(n4717), .B2(n4688), .ZN(n3634)
         );
  inv0d0 U5027 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[2]), .ZN(
        n5741) );
  oai22d1 U5028 ( .A1(n4718), .A2(n5741), .B1(n4717), .B2(n4689), .ZN(n3633)
         );
  inv0d0 U5029 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[3]), .ZN(
        n5742) );
  oai22d1 U5030 ( .A1(n4718), .A2(n5742), .B1(n4717), .B2(n4690), .ZN(n3632)
         );
  inv0d0 U5031 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[4]), .ZN(
        n5743) );
  oai22d1 U5032 ( .A1(n4718), .A2(n5743), .B1(n4717), .B2(n4691), .ZN(n3631)
         );
  inv0d0 U5033 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[5]), .ZN(
        n5744) );
  oai22d1 U5034 ( .A1(n4722), .A2(n5744), .B1(n4717), .B2(n4692), .ZN(n3630)
         );
  inv0d0 U5035 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[6]), .ZN(
        n5745) );
  oai22d1 U5036 ( .A1(n4722), .A2(n5745), .B1(n4717), .B2(n4693), .ZN(n3629)
         );
  inv0d0 U5037 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[7]), .ZN(
        n5746) );
  oai22d1 U5038 ( .A1(n4718), .A2(n5746), .B1(n4721), .B2(n4694), .ZN(n3628)
         );
  inv0d0 U5039 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[8]), .ZN(
        n5747) );
  oai22d1 U5040 ( .A1(n4722), .A2(n5747), .B1(n4717), .B2(n4695), .ZN(n3627)
         );
  inv0d0 U5041 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[9]), .ZN(
        n5748) );
  oai22d1 U5042 ( .A1(n4722), .A2(n5748), .B1(n4721), .B2(n4696), .ZN(n3626)
         );
  inv0d0 U5043 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[10]), .ZN(
        n5749) );
  oai22d1 U5044 ( .A1(n4722), .A2(n5749), .B1(n4717), .B2(n4697), .ZN(n3625)
         );
  inv0d0 U5045 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[11]), .ZN(
        n5750) );
  oai22d1 U5046 ( .A1(n4722), .A2(n5750), .B1(n4721), .B2(n4698), .ZN(n3624)
         );
  inv0d0 U5047 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[12]), .ZN(
        n5751) );
  oai22d1 U5048 ( .A1(n4722), .A2(n5751), .B1(n4717), .B2(n4699), .ZN(n3623)
         );
  inv0d0 U5049 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[13]), .ZN(
        n5752) );
  oai22d1 U5050 ( .A1(n4722), .A2(n5752), .B1(n4721), .B2(n4700), .ZN(n3622)
         );
  inv0d0 U5051 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[14]), .ZN(
        n5753) );
  oai22d1 U5052 ( .A1(n4718), .A2(n5753), .B1(n4721), .B2(n4701), .ZN(n3621)
         );
  inv0d0 U5053 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[15]), .ZN(
        n5754) );
  oai22d1 U5054 ( .A1(n4718), .A2(n5754), .B1(n4721), .B2(n4702), .ZN(n3620)
         );
  inv0d0 U5055 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[16]), .ZN(
        n5755) );
  oai22d1 U5056 ( .A1(n4722), .A2(n5755), .B1(n4717), .B2(n4703), .ZN(n3619)
         );
  inv0d0 U5057 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[17]), .ZN(
        n5756) );
  oai22d1 U5058 ( .A1(n4718), .A2(n5756), .B1(n4721), .B2(n4704), .ZN(n3618)
         );
  inv0d0 U5059 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[18]), .ZN(
        n5757) );
  oai22d1 U5060 ( .A1(n4718), .A2(n5757), .B1(n4721), .B2(n4705), .ZN(n3617)
         );
  inv0d0 U5061 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[19]), .ZN(
        n5758) );
  oai22d1 U5062 ( .A1(n4718), .A2(n5758), .B1(n4721), .B2(n4706), .ZN(n3616)
         );
  inv0d0 U5063 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[20]), .ZN(
        n5759) );
  oai22d1 U5064 ( .A1(n4718), .A2(n5759), .B1(n4721), .B2(n4707), .ZN(n3615)
         );
  inv0d0 U5065 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[21]), .ZN(
        n5760) );
  oai22d1 U5066 ( .A1(n4718), .A2(n5760), .B1(n4721), .B2(n4708), .ZN(n3614)
         );
  inv0d0 U5067 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[22]), .ZN(
        n5761) );
  oai22d1 U5068 ( .A1(n4718), .A2(n5761), .B1(n4721), .B2(n4709), .ZN(n3613)
         );
  inv0d0 U5069 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[23]), .ZN(
        n5762) );
  oai22d1 U5070 ( .A1(n4718), .A2(n5762), .B1(n4717), .B2(n4710), .ZN(n3612)
         );
  inv0d0 U5071 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[24]), .ZN(
        n5763) );
  oai22d1 U5072 ( .A1(n4722), .A2(n5763), .B1(n4717), .B2(n4711), .ZN(n3611)
         );
  inv0d0 U5073 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[25]), .ZN(
        n5764) );
  oai22d1 U5074 ( .A1(n4722), .A2(n5764), .B1(n4717), .B2(n4712), .ZN(n3610)
         );
  inv0d0 U5075 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[26]), .ZN(
        n5766) );
  oai22d1 U5076 ( .A1(n4722), .A2(n5766), .B1(n4717), .B2(n4713), .ZN(n3609)
         );
  inv0d0 U5077 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[27]), .ZN(
        n5769) );
  oai22d1 U5078 ( .A1(n4718), .A2(n5769), .B1(n4721), .B2(n4714), .ZN(n3608)
         );
  inv0d0 U5079 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[28]), .ZN(
        n5767) );
  oai22d1 U5080 ( .A1(n4722), .A2(n5767), .B1(n4721), .B2(n4715), .ZN(n3607)
         );
  inv0d0 U5081 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[29]), .ZN(
        n5773) );
  oai22d1 U5082 ( .A1(n4718), .A2(n5773), .B1(n4717), .B2(n4716), .ZN(n3606)
         );
  inv0d0 U5083 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[30]), .ZN(
        n5771) );
  oai22d1 U5084 ( .A1(n4722), .A2(n5771), .B1(n4721), .B2(n4719), .ZN(n3605)
         );
  inv0d0 U5085 ( .I(mgmtsoc_litespisdrphycore_source_payload_data[31]), .ZN(
        n5775) );
  oai22d1 U5086 ( .A1(n4722), .A2(n5775), .B1(n4721), .B2(n4720), .ZN(n3604)
         );
  or02d1 U5087 ( .A1(n4724), .A2(n5111), .Z(n4771) );
  oai21d1 U5088 ( .B1(n4957), .B2(n4723), .A(n4771), .ZN(n3603) );
  nd02d1 U5089 ( .A1(n5955), .A2(n4724), .ZN(n4760) );
  buffd1 U5090 ( .I(n4760), .Z(n4762) );
  buffd3 U5091 ( .I(n4771), .Z(n4767) );
  oai22d1 U5092 ( .A1(n5290), .A2(n4762), .B1(n4725), .B2(n4767), .ZN(n3602)
         );
  buffd1 U5093 ( .I(n4760), .Z(n4772) );
  oai22d1 U5094 ( .A1(n5294), .A2(n4772), .B1(n4726), .B2(n4767), .ZN(n3601)
         );
  oai22d1 U5095 ( .A1(n5245), .A2(n4772), .B1(n4727), .B2(n4767), .ZN(n3600)
         );
  inv0d0 U5096 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[3]), .ZN(
        n4728) );
  oai22d1 U5097 ( .A1(n5006), .A2(n4772), .B1(n4728), .B2(n4767), .ZN(n3599)
         );
  inv0d0 U5098 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[4]), .ZN(
        n4729) );
  oai22d1 U5099 ( .A1(n5008), .A2(n4760), .B1(n4729), .B2(n4767), .ZN(n3598)
         );
  inv0d0 U5100 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[5]), .ZN(
        n4730) );
  oai22d1 U5101 ( .A1(n5010), .A2(n4772), .B1(n4730), .B2(n4767), .ZN(n3597)
         );
  inv0d0 U5102 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[6]), .ZN(
        n4731) );
  oai22d1 U5103 ( .A1(n5012), .A2(n4772), .B1(n4731), .B2(n4767), .ZN(n3596)
         );
  inv0d0 U5104 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[7]), .ZN(
        n4732) );
  oai22d1 U5105 ( .A1(n5251), .A2(n4762), .B1(n4732), .B2(n4767), .ZN(n3595)
         );
  inv0d0 U5106 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[8]), .ZN(
        n4733) );
  oai22d1 U5107 ( .A1(n4783), .A2(n4760), .B1(n4733), .B2(n4767), .ZN(n3594)
         );
  inv0d0 U5108 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[9]), .ZN(
        n4734) );
  oai22d1 U5109 ( .A1(n4593), .A2(n4762), .B1(n4734), .B2(n4767), .ZN(n3593)
         );
  inv0d0 U5110 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[10]), .ZN(
        n4735) );
  oai22d1 U5111 ( .A1(n4595), .A2(n4762), .B1(n4735), .B2(n4767), .ZN(n3592)
         );
  inv0d0 U5112 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[11]), .ZN(
        n4736) );
  oai22d1 U5113 ( .A1(n5254), .A2(n4762), .B1(n4736), .B2(n4767), .ZN(n3591)
         );
  inv0d0 U5114 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[12]), .ZN(
        n4737) );
  oai22d1 U5115 ( .A1(n4598), .A2(n4762), .B1(n4737), .B2(n4767), .ZN(n3590)
         );
  inv0d0 U5116 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[13]), .ZN(
        n4738) );
  oai22d1 U5117 ( .A1(n4790), .A2(n4762), .B1(n4738), .B2(n4767), .ZN(n3589)
         );
  inv0d0 U5118 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[14]), .ZN(
        n4739) );
  oai22d1 U5119 ( .A1(n4601), .A2(n4762), .B1(n4739), .B2(n4767), .ZN(n3588)
         );
  inv0d0 U5120 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[15]), .ZN(
        n4740) );
  oai22d1 U5121 ( .A1(n4793), .A2(n4762), .B1(n4740), .B2(n4767), .ZN(n3587)
         );
  inv0d0 U5122 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[16]), .ZN(
        n4741) );
  oai22d1 U5123 ( .A1(n2003), .A2(n4762), .B1(n4741), .B2(n4767), .ZN(n3586)
         );
  inv0d0 U5124 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[17]), .ZN(
        n4742) );
  oai22d1 U5125 ( .A1(n5259), .A2(n4762), .B1(n4742), .B2(n4767), .ZN(n3585)
         );
  inv0d0 U5126 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[18]), .ZN(
        n4743) );
  oai22d1 U5127 ( .A1(n5260), .A2(n4772), .B1(n4743), .B2(n4767), .ZN(n3584)
         );
  inv0d0 U5128 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[19]), .ZN(
        n4744) );
  oai22d1 U5129 ( .A1(n5262), .A2(n4760), .B1(n4744), .B2(n4767), .ZN(n3583)
         );
  inv0d0 U5130 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[20]), .ZN(
        n4745) );
  oai22d1 U5131 ( .A1(n5263), .A2(n4762), .B1(n4745), .B2(n4767), .ZN(n3582)
         );
  inv0d0 U5132 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[21]), .ZN(
        n4746) );
  oai22d1 U5133 ( .A1(n5264), .A2(n4760), .B1(n4746), .B2(n4767), .ZN(n3581)
         );
  inv0d0 U5134 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[22]), .ZN(
        n4747) );
  oai22d1 U5135 ( .A1(n5266), .A2(n4762), .B1(n4747), .B2(n4767), .ZN(n3580)
         );
  inv0d0 U5136 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[23]), .ZN(
        n4748) );
  oai22d1 U5137 ( .A1(n5268), .A2(n4772), .B1(n4748), .B2(n4767), .ZN(n3579)
         );
  inv0d0 U5138 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[24]), .ZN(
        n4749) );
  oai22d1 U5139 ( .A1(n5270), .A2(n4772), .B1(n4749), .B2(n4767), .ZN(n3578)
         );
  inv0d0 U5140 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[25]), .ZN(
        n4750) );
  oai22d1 U5141 ( .A1(n5271), .A2(n4762), .B1(n4750), .B2(n4767), .ZN(n3577)
         );
  inv0d0 U5142 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[26]), .ZN(
        n4751) );
  oai22d1 U5143 ( .A1(n5273), .A2(n4762), .B1(n4751), .B2(n4771), .ZN(n3576)
         );
  inv0d0 U5144 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[27]), .ZN(
        n4752) );
  oai22d1 U5145 ( .A1(n5275), .A2(n4760), .B1(n4752), .B2(n4771), .ZN(n3575)
         );
  inv0d0 U5146 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[28]), .ZN(
        n4753) );
  oai22d1 U5147 ( .A1(n5276), .A2(n4760), .B1(n4753), .B2(n4767), .ZN(n3574)
         );
  inv0d0 U5148 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[29]), .ZN(
        n4754) );
  oai22d1 U5149 ( .A1(n5280), .A2(n4760), .B1(n4754), .B2(n4771), .ZN(n3573)
         );
  inv0d0 U5150 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[30]), .ZN(
        n4755) );
  oai22d1 U5151 ( .A1(n5283), .A2(n4760), .B1(n4755), .B2(n4771), .ZN(n3572)
         );
  inv0d0 U5152 ( .I(mgmtsoc_port_master_user_port_sink_payload_data[31]), .ZN(
        n4756) );
  oai22d1 U5153 ( .A1(n5287), .A2(n4772), .B1(n4756), .B2(n4771), .ZN(n3571)
         );
  oai22d1 U5154 ( .A1(n4774), .A2(n4772), .B1(n4757), .B2(n4767), .ZN(n3570)
         );
  inv0d0 U5155 ( .I(mgmtsoc_master_tx_fifo_sink_payload_len[1]), .ZN(n4775) );
  inv0d0 U5156 ( .I(mgmtsoc_port_master_user_port_sink_payload_len[1]), .ZN(
        n4758) );
  oai22d1 U5157 ( .A1(n4775), .A2(n4762), .B1(n4758), .B2(n4771), .ZN(n3569)
         );
  inv0d0 U5158 ( .I(mgmtsoc_port_master_user_port_sink_payload_len[2]), .ZN(
        n4759) );
  oai22d1 U5159 ( .A1(n4776), .A2(n4760), .B1(n4759), .B2(n4767), .ZN(n3568)
         );
  inv0d0 U5160 ( .I(mgmtsoc_port_master_user_port_sink_payload_len[3]), .ZN(
        n4761) );
  oai22d1 U5161 ( .A1(n4777), .A2(n4762), .B1(n4761), .B2(n4767), .ZN(n3567)
         );
  inv0d0 U5162 ( .I(mgmtsoc_port_master_user_port_sink_payload_len[4]), .ZN(
        n4763) );
  oai22d1 U5163 ( .A1(n4778), .A2(n4772), .B1(n4763), .B2(n4771), .ZN(n3566)
         );
  oai22d1 U5164 ( .A1(n4779), .A2(n4772), .B1(n4764), .B2(n4771), .ZN(n3565)
         );
  oai22d1 U5165 ( .A1(n4782), .A2(n4772), .B1(n4765), .B2(n4767), .ZN(n3564)
         );
  oai22d1 U5166 ( .A1(n4784), .A2(n4772), .B1(n4766), .B2(n4767), .ZN(n3563)
         );
  oai22d1 U5167 ( .A1(n4785), .A2(n4772), .B1(n4768), .B2(n4767), .ZN(n3562)
         );
  oai22d1 U5168 ( .A1(n4786), .A2(n4772), .B1(n4769), .B2(n4771), .ZN(n3561)
         );
  inv0d0 U5169 ( .I(\mgmtsoc_port_master_user_port_sink_payload_mask[0] ), 
        .ZN(n4770) );
  oai22d1 U5170 ( .A1(n4794), .A2(n4772), .B1(n4771), .B2(n4770), .ZN(n3560)
         );
  buffd1 U5171 ( .I(n4795), .Z(n4805) );
  buffd1 U5172 ( .I(n4797), .Z(n4804) );
  oai22d1 U5173 ( .A1(n4808), .A2(n4805), .B1(n4804), .B2(n4774), .ZN(n3559)
         );
  oai22d1 U5174 ( .A1(n5294), .A2(n4805), .B1(n4804), .B2(n4775), .ZN(n3558)
         );
  oai22d1 U5175 ( .A1(n5245), .A2(n4805), .B1(n4804), .B2(n4776), .ZN(n3557)
         );
  oai22d1 U5176 ( .A1(n5006), .A2(n4805), .B1(n4797), .B2(n4777), .ZN(n3556)
         );
  oai22d1 U5177 ( .A1(n5008), .A2(n4805), .B1(n4804), .B2(n4778), .ZN(n3555)
         );
  oai22d1 U5178 ( .A1(n5010), .A2(n4805), .B1(n4797), .B2(n4779), .ZN(n3554)
         );
  oai22d1 U5179 ( .A1(n5012), .A2(n4805), .B1(n4797), .B2(n4780), .ZN(n3553)
         );
  oai22d1 U5180 ( .A1(n5251), .A2(n4805), .B1(n4804), .B2(n4781), .ZN(n3552)
         );
  oai22d1 U5181 ( .A1(n4783), .A2(n4795), .B1(n4797), .B2(n4782), .ZN(n3551)
         );
  oai22d1 U5182 ( .A1(n4593), .A2(n4795), .B1(n4797), .B2(n4784), .ZN(n3550)
         );
  oai22d1 U5183 ( .A1(n4595), .A2(n4795), .B1(n4804), .B2(n4785), .ZN(n3549)
         );
  oai22d1 U5184 ( .A1(n4787), .A2(n4795), .B1(n4804), .B2(n4786), .ZN(n3548)
         );
  oai22d1 U5185 ( .A1(n4598), .A2(n4795), .B1(n4797), .B2(n4788), .ZN(n3547)
         );
  oai22d1 U5186 ( .A1(n4790), .A2(n4795), .B1(n4804), .B2(n4789), .ZN(n3546)
         );
  oai22d1 U5187 ( .A1(n4601), .A2(n4795), .B1(n4804), .B2(n4791), .ZN(n3545)
         );
  oai22d1 U5188 ( .A1(n4793), .A2(n4805), .B1(n4804), .B2(n4792), .ZN(n3544)
         );
  oai22d1 U5189 ( .A1(n2003), .A2(n4795), .B1(n4797), .B2(n4794), .ZN(n3543)
         );
  oai22d1 U5190 ( .A1(n5259), .A2(n4805), .B1(n4797), .B2(n4796), .ZN(n3542)
         );
  oai22d1 U5191 ( .A1(n5260), .A2(n4805), .B1(n4804), .B2(n4798), .ZN(n3541)
         );
  oai22d1 U5192 ( .A1(n5262), .A2(n4805), .B1(n4804), .B2(n4799), .ZN(n3540)
         );
  oai22d1 U5193 ( .A1(n5263), .A2(n4805), .B1(n4804), .B2(n4800), .ZN(n3539)
         );
  oai22d1 U5194 ( .A1(n5264), .A2(n4805), .B1(n4804), .B2(n4801), .ZN(n3538)
         );
  oai22d1 U5195 ( .A1(n5266), .A2(n4805), .B1(n4804), .B2(n4802), .ZN(n3537)
         );
  oai22d1 U5196 ( .A1(n5268), .A2(n4805), .B1(n4804), .B2(n4803), .ZN(n3536)
         );
  an02d0 U5197 ( .A1(n4806), .A2(n5240), .Z(n4809) );
  oai21d1 U5198 ( .B1(\litespi_request[1] ), .B2(n4809), .A(n5319), .ZN(n4807)
         );
  aoi21d1 U5199 ( .B1(n4809), .B2(n5290), .A(n4807), .ZN(n3535) );
  oai21d1 U5200 ( .B1(n4811), .B2(n4810), .A(n5319), .ZN(n4819) );
  aoim22d1 U5201 ( .A1(n4955), .A2(n4819), .B1(
        mgmtsoc_litespimmap_spi_dummy_bits[0]), .B2(n4812), .Z(n3534) );
  inv0d0 U5202 ( .I(mgmtsoc_litespimmap_spi_dummy_bits[1]), .ZN(n4813) );
  oai22d1 U5203 ( .A1(n5294), .A2(n4821), .B1(n4813), .B2(n4819), .ZN(n3533)
         );
  oai22d1 U5204 ( .A1(n5004), .A2(n4821), .B1(n4814), .B2(n4819), .ZN(n3532)
         );
  oai22d1 U5205 ( .A1(n5006), .A2(n4821), .B1(n4815), .B2(n4819), .ZN(n3531)
         );
  oai22d1 U5206 ( .A1(n5008), .A2(n4821), .B1(n4816), .B2(n4819), .ZN(n3530)
         );
  oai22d1 U5207 ( .A1(n5010), .A2(n4821), .B1(n4817), .B2(n4819), .ZN(n3529)
         );
  oai22d1 U5208 ( .A1(n5012), .A2(n4821), .B1(n4818), .B2(n4819), .ZN(n3528)
         );
  oai22d1 U5209 ( .A1(n5251), .A2(n4821), .B1(n4820), .B2(n4819), .ZN(n3527)
         );
  nr04d0 U5210 ( .A1(mgmtsoc_litespimmap_count[3]), .A2(
        mgmtsoc_litespimmap_count[2]), .A3(mgmtsoc_litespimmap_count[1]), .A4(
        mgmtsoc_litespimmap_count[0]), .ZN(n4832) );
  inv0d0 U5211 ( .I(mgmtsoc_litespimmap_count[4]), .ZN(n4831) );
  nd02d0 U5212 ( .A1(n4832), .A2(n4831), .ZN(n4830) );
  nr02d0 U5213 ( .A1(mgmtsoc_litespimmap_count[5]), .A2(n4830), .ZN(n4828) );
  inv0d0 U5214 ( .I(mgmtsoc_litespimmap_count[6]), .ZN(n4827) );
  nd02d0 U5215 ( .A1(n4828), .A2(n4827), .ZN(n4826) );
  nr02d0 U5216 ( .A1(mgmtsoc_litespimmap_count[7]), .A2(n4826), .ZN(n4824) );
  inv0d0 U5217 ( .I(mgmtsoc_litespimmap_count[8]), .ZN(n4823) );
  nd02d0 U5218 ( .A1(n4824), .A2(n4823), .ZN(n4842) );
  nr02d0 U5219 ( .A1(mgmtsoc_litespimmap_count[0]), .A2(n4834), .ZN(n3526) );
  oai211d1 U5220 ( .C1(n4824), .C2(n4823), .A(n4822), .B(n4881), .ZN(n3525) );
  inv0d0 U5221 ( .I(n4834), .ZN(n4837) );
  aon211d1 U5222 ( .C1(mgmtsoc_litespimmap_count[7]), .C2(n4826), .B(n4824), 
        .A(n4837), .ZN(n4825) );
  inv0d0 U5223 ( .I(n4825), .ZN(n3524) );
  oan211d1 U5224 ( .C1(n4828), .C2(n4827), .B(n4826), .A(n4834), .ZN(n3523) );
  aon211d1 U5225 ( .C1(mgmtsoc_litespimmap_count[5]), .C2(n4830), .B(n4828), 
        .A(n4837), .ZN(n4829) );
  inv0d0 U5226 ( .I(n4829), .ZN(n3522) );
  oan211d1 U5227 ( .C1(n4832), .C2(n4831), .B(n4830), .A(n4834), .ZN(n3521) );
  or03d0 U5228 ( .A1(mgmtsoc_litespimmap_count[2]), .A2(
        mgmtsoc_litespimmap_count[1]), .A3(mgmtsoc_litespimmap_count[0]), .Z(
        n4835) );
  aon211d1 U5229 ( .C1(n4835), .C2(mgmtsoc_litespimmap_count[3]), .B(n4832), 
        .A(n4837), .ZN(n4833) );
  inv0d0 U5230 ( .I(n4833), .ZN(n3520) );
  nr02d0 U5231 ( .A1(mgmtsoc_litespimmap_count[1]), .A2(
        mgmtsoc_litespimmap_count[0]), .ZN(n4838) );
  inv0d0 U5232 ( .I(mgmtsoc_litespimmap_count[2]), .ZN(n4836) );
  oan211d1 U5233 ( .C1(n4838), .C2(n4836), .B(n4835), .A(n4834), .ZN(n3519) );
  aon211d1 U5234 ( .C1(mgmtsoc_litespimmap_count[1]), .C2(
        mgmtsoc_litespimmap_count[0]), .B(n4838), .A(n4837), .ZN(n4839) );
  inv0d0 U5235 ( .I(n4839), .ZN(n3518) );
  nd02d0 U5236 ( .A1(n4841), .A2(n4840), .ZN(n5729) );
  inv0d0 U5237 ( .I(n5729), .ZN(n5707) );
  inv0d2 U5238 ( .I(n5707), .ZN(n5721) );
  oai21d1 U5239 ( .B1(n4843), .B2(n4842), .A(mgmtsoc_litespimmap_burst_cs), 
        .ZN(n4844) );
  oan211d1 U5240 ( .C1(n4845), .C2(n5721), .B(n4844), .A(n4878), .ZN(n3517) );
  oan211d1 U5241 ( .C1(litespi_tx_mux_sel), .C2(n4847), .B(n4846), .A(sys_rst), 
        .ZN(n4853) );
  oai21d1 U5242 ( .B1(mgmtsoc_litespisdrphycore_count[0]), .B2(n4856), .A(
        n4853), .ZN(n3516) );
  nr03d0 U5243 ( .A1(mgmtsoc_litespisdrphycore_count[2]), .A2(
        mgmtsoc_litespisdrphycore_count[1]), .A3(
        mgmtsoc_litespisdrphycore_count[0]), .ZN(n4851) );
  inv0d0 U5244 ( .I(mgmtsoc_litespisdrphycore_count[3]), .ZN(n4848) );
  oai21d1 U5245 ( .B1(n4851), .B2(n4848), .A(n4853), .ZN(n3515) );
  oai21d1 U5246 ( .B1(mgmtsoc_litespisdrphycore_count[1]), .B2(
        mgmtsoc_litespisdrphycore_count[0]), .A(
        mgmtsoc_litespisdrphycore_count[2]), .ZN(n4849) );
  inv0d0 U5247 ( .I(n4849), .ZN(n4850) );
  aon211d1 U5248 ( .C1(mgmtsoc_litespisdrphycore_count[3]), .C2(n4851), .B(
        n4850), .A(n4853), .ZN(n4852) );
  inv0d0 U5249 ( .I(n4852), .ZN(n3514) );
  inv0d0 U5250 ( .I(mgmtsoc_litespisdrphycore_count[1]), .ZN(n4855) );
  inv0d0 U5251 ( .I(mgmtsoc_litespisdrphycore_count[0]), .ZN(n4854) );
  oai321d1 U5252 ( .C1(mgmtsoc_litespisdrphycore_count[1]), .C2(
        mgmtsoc_litespisdrphycore_count[0]), .C3(n4856), .B1(n4855), .B2(n4854), .A(n4853), .ZN(n3513) );
  oai211d1 U5253 ( .C1(n4859), .C2(mgmtsoc_litespisdrphycore_clk), .A(n4857), 
        .B(n5340), .ZN(n4858) );
  aoi21d1 U5254 ( .B1(n4859), .B2(mgmtsoc_litespisdrphycore_clk), .A(n4858), 
        .ZN(n3512) );
  inv0d0 U5255 ( .I(n4861), .ZN(n4870) );
  aoim22d1 U5256 ( .A1(n4861), .A2(n5290), .B1(n4871), .B2(
        mgmtsoc_litespisdrphycore_div[0]), .Z(n3511) );
  oai22d1 U5257 ( .A1(n4863), .A2(n4871), .B1(n4862), .B2(n4870), .ZN(n3510)
         );
  oai22d1 U5258 ( .A1(n4864), .A2(n4871), .B1(n5004), .B2(n4870), .ZN(n3509)
         );
  oai22d1 U5259 ( .A1(n4865), .A2(n4871), .B1(n5246), .B2(n4870), .ZN(n3508)
         );
  oai22d1 U5260 ( .A1(n4867), .A2(n4871), .B1(n4866), .B2(n4870), .ZN(n3507)
         );
  oai22d1 U5261 ( .A1(n4868), .A2(n4871), .B1(n5248), .B2(n4870), .ZN(n3506)
         );
  oai22d1 U5262 ( .A1(n4869), .A2(n4871), .B1(n5249), .B2(n4870), .ZN(n3505)
         );
  oai22d1 U5263 ( .A1(n4872), .A2(n4871), .B1(n5251), .B2(n4870), .ZN(n3504)
         );
  nd02d0 U5264 ( .A1(n4873), .A2(n4997), .ZN(n4875) );
  nd03d0 U5265 ( .A1(n4875), .A2(mgmtsoc_zero2), .A3(n5301), .ZN(n4874) );
  oai21d1 U5266 ( .B1(n4875), .B2(n4955), .A(n4874), .ZN(n3503) );
  oai21d1 U5267 ( .B1(n4877), .B2(n4955), .A(n4876), .ZN(n3502) );
  oaim21d1 U5268 ( .B1(mgmtsoc_pending_r), .B2(mgmtsoc_pending_re), .A(
        mgmtsoc_zero1), .ZN(n4879) );
  oan211d1 U5269 ( .C1(mgmtsoc_zero_trigger_d), .C2(n4880), .B(n4879), .A(
        n4878), .ZN(n3501) );
  inv0d0 U5270 ( .I(csrbank10_value_w[0]), .ZN(n4883) );
  or02d1 U5271 ( .A1(mgmtsoc_update_value_re), .A2(n5100), .Z(n4934) );
  nd02d1 U5272 ( .A1(mgmtsoc_update_value_re), .A2(n5956), .ZN(n4948) );
  oai22d1 U5273 ( .A1(n4883), .A2(n4934), .B1(n4882), .B2(n4948), .ZN(n3500)
         );
  inv0d0 U5274 ( .I(mgmtsoc_value[1]), .ZN(n4885) );
  buffd1 U5275 ( .I(n4948), .Z(n4944) );
  oai22d1 U5276 ( .A1(n4885), .A2(n4944), .B1(n4884), .B2(n4934), .ZN(n3499)
         );
  oai22d1 U5277 ( .A1(n4887), .A2(n4944), .B1(n4886), .B2(n4934), .ZN(n3498)
         );
  inv0d0 U5278 ( .I(mgmtsoc_value[3]), .ZN(n4889) );
  oai22d1 U5279 ( .A1(n4889), .A2(n4948), .B1(n4888), .B2(n4934), .ZN(n3497)
         );
  inv0d0 U5280 ( .I(mgmtsoc_value[4]), .ZN(n4891) );
  oai22d1 U5281 ( .A1(n4891), .A2(n4944), .B1(n4890), .B2(n4934), .ZN(n3496)
         );
  buffd1 U5282 ( .I(n4934), .Z(n4946) );
  oai22d1 U5283 ( .A1(n4893), .A2(n4944), .B1(n4892), .B2(n4946), .ZN(n3495)
         );
  inv0d0 U5284 ( .I(mgmtsoc_value[6]), .ZN(n4895) );
  oai22d1 U5285 ( .A1(n4895), .A2(n4944), .B1(n4894), .B2(n4934), .ZN(n3494)
         );
  oai22d1 U5286 ( .A1(n4897), .A2(n4944), .B1(n4896), .B2(n4934), .ZN(n3493)
         );
  inv0d0 U5287 ( .I(mgmtsoc_value[8]), .ZN(n4899) );
  oai22d1 U5288 ( .A1(n4899), .A2(n4944), .B1(n4898), .B2(n4934), .ZN(n3492)
         );
  inv0d0 U5289 ( .I(mgmtsoc_value[9]), .ZN(n4901) );
  oai22d1 U5290 ( .A1(n4901), .A2(n4944), .B1(n4900), .B2(n4946), .ZN(n3491)
         );
  inv0d0 U5291 ( .I(mgmtsoc_value[10]), .ZN(n4903) );
  oai22d1 U5292 ( .A1(n4903), .A2(n4944), .B1(n4902), .B2(n4946), .ZN(n3490)
         );
  oai22d1 U5293 ( .A1(n4905), .A2(n4944), .B1(n4904), .B2(n4946), .ZN(n3489)
         );
  inv0d0 U5294 ( .I(mgmtsoc_value[12]), .ZN(n4907) );
  oai22d1 U5295 ( .A1(n4907), .A2(n4944), .B1(n4906), .B2(n4946), .ZN(n3488)
         );
  oai22d1 U5296 ( .A1(n4909), .A2(n4944), .B1(n4908), .B2(n4946), .ZN(n3487)
         );
  inv0d0 U5297 ( .I(mgmtsoc_value[14]), .ZN(n4911) );
  oai22d1 U5298 ( .A1(n4911), .A2(n4944), .B1(n4910), .B2(n4946), .ZN(n3486)
         );
  oai22d1 U5299 ( .A1(n4913), .A2(n4948), .B1(n4912), .B2(n4946), .ZN(n3485)
         );
  inv0d0 U5300 ( .I(mgmtsoc_value[16]), .ZN(n4915) );
  oai22d1 U5301 ( .A1(n4915), .A2(n4944), .B1(n4914), .B2(n4946), .ZN(n3484)
         );
  oai22d1 U5302 ( .A1(n4917), .A2(n4948), .B1(n4916), .B2(n4946), .ZN(n3483)
         );
  inv0d0 U5303 ( .I(mgmtsoc_value[18]), .ZN(n4919) );
  oai22d1 U5304 ( .A1(n4919), .A2(n4944), .B1(n4918), .B2(n4946), .ZN(n3482)
         );
  oai22d1 U5305 ( .A1(n4921), .A2(n4944), .B1(n4920), .B2(n4934), .ZN(n3481)
         );
  inv0d0 U5306 ( .I(mgmtsoc_value[20]), .ZN(n4923) );
  oai22d1 U5307 ( .A1(n4923), .A2(n4948), .B1(n4922), .B2(n4934), .ZN(n3480)
         );
  oai22d1 U5308 ( .A1(n4925), .A2(n4948), .B1(n4924), .B2(n4934), .ZN(n3479)
         );
  inv0d0 U5309 ( .I(mgmtsoc_value[22]), .ZN(n4927) );
  oai22d1 U5310 ( .A1(n4927), .A2(n4948), .B1(n4926), .B2(n4934), .ZN(n3478)
         );
  oai22d1 U5311 ( .A1(n4929), .A2(n4948), .B1(n4928), .B2(n4934), .ZN(n3477)
         );
  inv0d0 U5312 ( .I(mgmtsoc_value[24]), .ZN(n4931) );
  oai22d1 U5313 ( .A1(n4931), .A2(n4948), .B1(n4930), .B2(n4934), .ZN(n3476)
         );
  oai22d1 U5314 ( .A1(n4933), .A2(n4948), .B1(n4932), .B2(n4946), .ZN(n3475)
         );
  inv0d0 U5315 ( .I(mgmtsoc_value[26]), .ZN(n4936) );
  oai22d1 U5316 ( .A1(n4936), .A2(n4948), .B1(n4935), .B2(n4934), .ZN(n3474)
         );
  oai22d1 U5317 ( .A1(n4938), .A2(n4948), .B1(n4937), .B2(n4946), .ZN(n3473)
         );
  inv0d0 U5318 ( .I(mgmtsoc_value[28]), .ZN(n4940) );
  oai22d1 U5319 ( .A1(n4940), .A2(n4948), .B1(n4939), .B2(n4946), .ZN(n3472)
         );
  oai22d1 U5320 ( .A1(n4942), .A2(n4948), .B1(n4941), .B2(n4946), .ZN(n3471)
         );
  inv0d0 U5321 ( .I(mgmtsoc_value[30]), .ZN(n4945) );
  oai22d1 U5322 ( .A1(n4945), .A2(n4944), .B1(n4943), .B2(n4946), .ZN(n3470)
         );
  inv0d0 U5323 ( .I(mgmtsoc_value[31]), .ZN(n4949) );
  oai22d1 U5324 ( .A1(n4949), .A2(n4948), .B1(n4947), .B2(n4946), .ZN(n3469)
         );
  oai21d1 U5325 ( .B1(n4951), .B2(n4955), .A(n4950), .ZN(n3468) );
  nd02d0 U5326 ( .A1(n4952), .A2(n4997), .ZN(n4953) );
  inv0d0 U5327 ( .I(n4953), .ZN(n4956) );
  aoi22d1 U5328 ( .A1(n4956), .A2(n4955), .B1(n4954), .B2(n4953), .ZN(n3467)
         );
  or02d1 U5329 ( .A1(n4958), .A2(n4957), .Z(n4996) );
  oai21d1 U5330 ( .B1(n4960), .B2(n4959), .A(n4881), .ZN(n4987) );
  oai22d1 U5331 ( .A1(n5290), .A2(n4996), .B1(n4961), .B2(n4987), .ZN(n3466)
         );
  buffd1 U5332 ( .I(n4987), .Z(n4994) );
  oai22d1 U5333 ( .A1(n5294), .A2(n4996), .B1(n4962), .B2(n4994), .ZN(n3465)
         );
  oai22d1 U5334 ( .A1(n5004), .A2(n4996), .B1(n4963), .B2(n4987), .ZN(n3464)
         );
  buffd1 U5335 ( .I(n4996), .Z(n4991) );
  oai22d1 U5336 ( .A1(n5006), .A2(n4991), .B1(n4964), .B2(n4994), .ZN(n3463)
         );
  oai22d1 U5337 ( .A1(n5008), .A2(n4991), .B1(n4965), .B2(n4994), .ZN(n3462)
         );
  oai22d1 U5338 ( .A1(n5010), .A2(n4991), .B1(n4966), .B2(n4994), .ZN(n3461)
         );
  oai22d1 U5339 ( .A1(n5012), .A2(n4996), .B1(n4967), .B2(n4994), .ZN(n3460)
         );
  oai22d1 U5340 ( .A1(n5251), .A2(n4996), .B1(n4968), .B2(n4994), .ZN(n3459)
         );
  oai22d1 U5341 ( .A1(n5015), .A2(n4991), .B1(n4969), .B2(n4994), .ZN(n3458)
         );
  oai22d1 U5342 ( .A1(n5017), .A2(n4991), .B1(n4970), .B2(n4994), .ZN(n3457)
         );
  oai22d1 U5343 ( .A1(n5019), .A2(n4991), .B1(n4971), .B2(n4987), .ZN(n3456)
         );
  oai22d1 U5344 ( .A1(n4787), .A2(n4991), .B1(n4972), .B2(n4987), .ZN(n3455)
         );
  oai22d1 U5345 ( .A1(n5022), .A2(n4991), .B1(n4973), .B2(n4994), .ZN(n3454)
         );
  oai22d1 U5346 ( .A1(n5024), .A2(n4991), .B1(n4974), .B2(n4987), .ZN(n3453)
         );
  oai22d1 U5347 ( .A1(n5026), .A2(n4991), .B1(n4975), .B2(n4987), .ZN(n3452)
         );
  oai22d1 U5348 ( .A1(n5028), .A2(n4991), .B1(n4976), .B2(n4987), .ZN(n3451)
         );
  oai22d1 U5349 ( .A1(n2003), .A2(n4991), .B1(n4977), .B2(n4987), .ZN(n3450)
         );
  oai22d1 U5350 ( .A1(n5259), .A2(n4991), .B1(n4978), .B2(n4987), .ZN(n3449)
         );
  oai22d1 U5351 ( .A1(n5260), .A2(n4996), .B1(n4979), .B2(n4987), .ZN(n3448)
         );
  oai22d1 U5352 ( .A1(n5262), .A2(n4996), .B1(n4980), .B2(n4994), .ZN(n3447)
         );
  oai22d1 U5353 ( .A1(n5263), .A2(n4991), .B1(n4981), .B2(n4987), .ZN(n3446)
         );
  oai22d1 U5354 ( .A1(n5264), .A2(n4996), .B1(n4982), .B2(n4994), .ZN(n3445)
         );
  oai22d1 U5355 ( .A1(n5266), .A2(n4996), .B1(n4983), .B2(n4987), .ZN(n3444)
         );
  oai22d1 U5356 ( .A1(n5268), .A2(n4996), .B1(n4984), .B2(n4994), .ZN(n3443)
         );
  oai22d1 U5357 ( .A1(n5270), .A2(n4996), .B1(n4985), .B2(n4987), .ZN(n3442)
         );
  oai22d1 U5358 ( .A1(n5271), .A2(n4996), .B1(n4986), .B2(n4987), .ZN(n3441)
         );
  oai22d1 U5359 ( .A1(n5273), .A2(n4991), .B1(n4988), .B2(n4987), .ZN(n3440)
         );
  oai22d1 U5360 ( .A1(n5275), .A2(n4991), .B1(n4989), .B2(n4994), .ZN(n3439)
         );
  oai22d1 U5361 ( .A1(n5276), .A2(n4991), .B1(n4990), .B2(n4994), .ZN(n3438)
         );
  oai22d1 U5362 ( .A1(n5280), .A2(n4996), .B1(n4992), .B2(n4994), .ZN(n3437)
         );
  oai22d1 U5363 ( .A1(n5283), .A2(n4996), .B1(n4993), .B2(n4994), .ZN(n3436)
         );
  oai22d1 U5364 ( .A1(n5287), .A2(n4996), .B1(n4995), .B2(n4994), .ZN(n3435)
         );
  nd02d1 U5365 ( .A1(n5288), .A2(n5001), .ZN(n5038) );
  aoi22d1 U5366 ( .A1(n5000), .A2(n5038), .B1(n4999), .B2(n5001), .ZN(n3434)
         );
  nd12d1 U5367 ( .A1(n5001), .A2(n5340), .ZN(n5048) );
  buffd1 U5368 ( .I(n5048), .Z(n5045) );
  buffd1 U5369 ( .I(n5038), .Z(n5046) );
  oai22d1 U5370 ( .A1(n5294), .A2(n5045), .B1(n5002), .B2(n5046), .ZN(n3433)
         );
  oai22d1 U5371 ( .A1(n5004), .A2(n5045), .B1(n5003), .B2(n5038), .ZN(n3432)
         );
  oai22d1 U5372 ( .A1(n5006), .A2(n5045), .B1(n5005), .B2(n5046), .ZN(n3431)
         );
  oai22d1 U5373 ( .A1(n5008), .A2(n5045), .B1(n5007), .B2(n5038), .ZN(n3430)
         );
  oai22d1 U5374 ( .A1(n5010), .A2(n5045), .B1(n5009), .B2(n5046), .ZN(n3429)
         );
  oai22d1 U5375 ( .A1(n5012), .A2(n5045), .B1(n5011), .B2(n5038), .ZN(n3428)
         );
  oai22d1 U5376 ( .A1(n5251), .A2(n5045), .B1(n5013), .B2(n5046), .ZN(n3427)
         );
  oai22d1 U5377 ( .A1(n5015), .A2(n5045), .B1(n5014), .B2(n5038), .ZN(n3426)
         );
  oai22d1 U5378 ( .A1(n5017), .A2(n5045), .B1(n5016), .B2(n5046), .ZN(n3425)
         );
  oai22d1 U5379 ( .A1(n5019), .A2(n5045), .B1(n5018), .B2(n5038), .ZN(n3424)
         );
  oai22d1 U5380 ( .A1(n4787), .A2(n5048), .B1(n5020), .B2(n5038), .ZN(n3423)
         );
  oai22d1 U5381 ( .A1(n5022), .A2(n5048), .B1(n5021), .B2(n5038), .ZN(n3422)
         );
  oai22d1 U5382 ( .A1(n5024), .A2(n5048), .B1(n5023), .B2(n5038), .ZN(n3421)
         );
  oai22d1 U5383 ( .A1(n5026), .A2(n5045), .B1(n5025), .B2(n5038), .ZN(n3420)
         );
  oai22d1 U5384 ( .A1(n5028), .A2(n5048), .B1(n5027), .B2(n5038), .ZN(n3419)
         );
  oai22d1 U5385 ( .A1(n2003), .A2(n5045), .B1(n5029), .B2(n5046), .ZN(n3418)
         );
  oai22d1 U5386 ( .A1(n5259), .A2(n5048), .B1(n5030), .B2(n5046), .ZN(n3417)
         );
  oai22d1 U5387 ( .A1(n5260), .A2(n5045), .B1(n5031), .B2(n5038), .ZN(n3416)
         );
  oai22d1 U5388 ( .A1(n5262), .A2(n5048), .B1(n5032), .B2(n5046), .ZN(n3415)
         );
  oai22d1 U5389 ( .A1(n5263), .A2(n5048), .B1(n5033), .B2(n5046), .ZN(n3414)
         );
  oai22d1 U5390 ( .A1(n5264), .A2(n5048), .B1(n5034), .B2(n5038), .ZN(n3413)
         );
  oai22d1 U5391 ( .A1(n5266), .A2(n5048), .B1(n5035), .B2(n5038), .ZN(n3412)
         );
  oai22d1 U5392 ( .A1(n5268), .A2(n5048), .B1(n5036), .B2(n5046), .ZN(n3411)
         );
  oai22d1 U5393 ( .A1(n5270), .A2(n5045), .B1(n5037), .B2(n5046), .ZN(n3410)
         );
  oai22d1 U5394 ( .A1(n5271), .A2(n5045), .B1(n5039), .B2(n5038), .ZN(n3409)
         );
  oai22d1 U5395 ( .A1(n5273), .A2(n5048), .B1(n5040), .B2(n5046), .ZN(n3408)
         );
  oai22d1 U5396 ( .A1(n5275), .A2(n5048), .B1(n5041), .B2(n5046), .ZN(n3407)
         );
  oai22d1 U5397 ( .A1(n5276), .A2(n5045), .B1(n5042), .B2(n5046), .ZN(n3406)
         );
  oai22d1 U5398 ( .A1(n5280), .A2(n5048), .B1(n5043), .B2(n5046), .ZN(n3405)
         );
  oai22d1 U5399 ( .A1(n5283), .A2(n5045), .B1(n5044), .B2(n5046), .ZN(n3404)
         );
  oai22d1 U5400 ( .A1(n5287), .A2(n5048), .B1(n5047), .B2(n5046), .ZN(n3403)
         );
  nr02d0 U5401 ( .A1(mgmtsoc_vexriscv_i_cmd_valid), .A2(n5051), .ZN(n5055) );
  inv0d0 U5402 ( .I(mgmtsoc_vexriscv_i_cmd_valid), .ZN(n5099) );
  inv0d0 U5403 ( .I(mgmtsoc_vexriscv_transfer_complete), .ZN(n5056) );
  inv0d0 U5404 ( .I(mgmtsoc_vexriscv_transfer_wait_for_ack), .ZN(n5054) );
  an02d0 U5405 ( .A1(n5288), .A2(n5057), .Z(n5089) );
  buffd1 U5406 ( .I(n5089), .Z(n5085) );
  nd02d0 U5407 ( .A1(mgmtsoc_vexriscv_debug_bus_ack), .A2(n5085), .ZN(n5052)
         );
  nd03d0 U5408 ( .A1(mgmtsoc_vexriscv_transfer_complete), .A2(n5956), .A3(
        n5099), .ZN(n5053) );
  aon211d1 U5409 ( .C1(mgmtsoc_vexriscv_transfer_wait_for_ack), .C2(n5055), 
        .B(n5052), .A(n5053), .ZN(n3402) );
  oai31d1 U5410 ( .B1(n4878), .B2(n5055), .B3(n5054), .A(n5053), .ZN(n3401) );
  inv0d0 U5411 ( .I(mgmtsoc_vexriscv_o_cmd_ready), .ZN(n5095) );
  aoi211d1 U5412 ( .C1(n5056), .C2(n5095), .A(n4878), .B(n5099), .ZN(n3400) );
  nd12d0 U5413 ( .A1(n5057), .A2(n5956), .ZN(n5077) );
  buffd1 U5414 ( .I(n5077), .Z(n5093) );
  oaim22d1 U5415 ( .A1(n5058), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[0]), .B2(n5085), .ZN(n3399) );
  oaim22d1 U5416 ( .A1(n5059), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[1]), .B2(n5085), .ZN(n3398) );
  buffd1 U5417 ( .I(n5077), .Z(n5098) );
  oaim22d1 U5418 ( .A1(n5060), .A2(n5098), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[2]), .B2(n5085), .ZN(n3397) );
  oaim22d1 U5419 ( .A1(n5061), .A2(n5077), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[3]), .B2(n5085), .ZN(n3396) );
  oaim22d1 U5420 ( .A1(n5062), .A2(n5077), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[4]), .B2(n5085), .ZN(n3395) );
  buffd1 U5421 ( .I(n5089), .Z(n5094) );
  oaim22d1 U5422 ( .A1(n5063), .A2(n5098), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[5]), .B2(n5094), .ZN(n3394) );
  oaim22d1 U5423 ( .A1(n5064), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[6]), .B2(n5085), .ZN(n3393) );
  oaim22d1 U5424 ( .A1(n5065), .A2(n5098), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[7]), .B2(n5089), .ZN(n3392) );
  oaim22d1 U5425 ( .A1(n5066), .A2(n5077), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[8]), .B2(n5094), .ZN(n3391) );
  oaim22d1 U5426 ( .A1(n5067), .A2(n5098), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[9]), .B2(n5085), .ZN(n3390) );
  oaim22d1 U5427 ( .A1(n5068), .A2(n5098), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[10]), .B2(n5094), .ZN(n3389) );
  oaim22d1 U5428 ( .A1(n5069), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[11]), .B2(n5094), .ZN(n3388) );
  oaim22d1 U5429 ( .A1(n5070), .A2(n5077), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[12]), .B2(n5094), .ZN(n3387) );
  oaim22d1 U5430 ( .A1(n5071), .A2(n5098), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[13]), .B2(n5085), .ZN(n3386) );
  oaim22d1 U5431 ( .A1(n5072), .A2(n5098), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[14]), .B2(n5085), .ZN(n3385) );
  oaim22d1 U5432 ( .A1(n5073), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[15]), .B2(n5085), .ZN(n3384) );
  oaim22d1 U5433 ( .A1(n5074), .A2(n5077), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[16]), .B2(n5094), .ZN(n3383) );
  oaim22d1 U5434 ( .A1(n5075), .A2(n5098), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[17]), .B2(n5085), .ZN(n3382) );
  oaim22d1 U5435 ( .A1(n5076), .A2(n5098), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[18]), .B2(n5085), .ZN(n3381) );
  oaim22d1 U5436 ( .A1(n5078), .A2(n5077), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[19]), .B2(n5085), .ZN(n3380) );
  oaim22d1 U5437 ( .A1(n5079), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[20]), .B2(n5094), .ZN(n3379) );
  oaim22d1 U5438 ( .A1(n5080), .A2(n5098), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[21]), .B2(n5085), .ZN(n3378) );
  oaim22d1 U5439 ( .A1(n5081), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[22]), .B2(n5089), .ZN(n3377) );
  oaim22d1 U5440 ( .A1(n5082), .A2(n5098), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[23]), .B2(n5089), .ZN(n3376) );
  oaim22d1 U5441 ( .A1(n5083), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[24]), .B2(n5089), .ZN(n3375) );
  oaim22d1 U5442 ( .A1(n5084), .A2(n5098), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[25]), .B2(n5089), .ZN(n3374) );
  oaim22d1 U5443 ( .A1(n5086), .A2(n5098), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[26]), .B2(n5085), .ZN(n3373) );
  oaim22d1 U5444 ( .A1(n5087), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[27]), .B2(n5094), .ZN(n3372) );
  oaim22d1 U5445 ( .A1(n5088), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[28]), .B2(n5089), .ZN(n3371) );
  oaim22d1 U5446 ( .A1(n5090), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[29]), .B2(n5089), .ZN(n3370) );
  oaim22d1 U5447 ( .A1(n5091), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[30]), .B2(n5094), .ZN(n3369) );
  oaim22d1 U5448 ( .A1(n5092), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_data[31]), .B2(n5094), .ZN(n3368) );
  oaim22d1 U5449 ( .A1(n5611), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_address[2]), .B2(n5094), .ZN(n3367) );
  oaim22d1 U5450 ( .A1(n5614), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_address[3]), .B2(n5094), .ZN(n3366) );
  oaim22d1 U5451 ( .A1(n5617), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_address[4]), .B2(n5094), .ZN(n3365) );
  oaim22d1 U5452 ( .A1(n5621), .A2(n5093), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_address[5]), .B2(n5094), .ZN(n3364) );
  oaim22d1 U5453 ( .A1(n5625), .A2(n5098), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_address[6]), .B2(n5094), .ZN(n3363) );
  oaim22d1 U5454 ( .A1(n5629), .A2(n5098), .B1(
        mgmtsoc_vexriscv_i_cmd_payload_address[7]), .B2(n5094), .ZN(n3362) );
  oai211d1 U5455 ( .C1(n5099), .C2(n5095), .A(n5094), .B(
        mgmtsoc_vexriscv_i_cmd_payload_wr), .ZN(n5096) );
  oai21d1 U5456 ( .B1(n5097), .B2(n5098), .A(n5096), .ZN(n3361) );
  oai31d1 U5457 ( .B1(n5100), .B2(mgmtsoc_vexriscv_o_cmd_ready), .B3(n5099), 
        .A(n5098), .ZN(n3360) );
  nr04d0 U5458 ( .A1(n5156), .A2(n5152), .A3(n5148), .A4(n5144), .ZN(n5104) );
  nr04d0 U5459 ( .A1(n5113), .A2(n5124), .A3(n5120), .A4(n5116), .ZN(n5102) );
  nr04d0 U5460 ( .A1(n5140), .A2(n5136), .A3(n5132), .A4(n5128), .ZN(n5101) );
  nr04d0 U5461 ( .A1(n5222), .A2(n5218), .A3(n5213), .A4(n5209), .ZN(n5108) );
  nr04d0 U5462 ( .A1(n5239), .A2(n5234), .A3(n5230), .A4(n5226), .ZN(n5107) );
  nr04d0 U5463 ( .A1(n5188), .A2(n5184), .A3(n5180), .A4(n5176), .ZN(n5106) );
  nr04d0 U5464 ( .A1(n5205), .A2(n5200), .A3(n5196), .A4(n5192), .ZN(n5105) );
  oai21d1 U5465 ( .B1(n5110), .B2(n5109), .A(n5335), .ZN(n5112) );
  nd02d1 U5466 ( .A1(n5288), .A2(n5112), .ZN(n5204) );
  or02d1 U5467 ( .A1(n5112), .A2(n5111), .Z(n5217) );
  aoi22d1 U5468 ( .A1(mgmtsoc_bus_errors_status[0]), .A2(n5204), .B1(n5217), 
        .B2(n5113), .ZN(n3359) );
  xn02d1 U5469 ( .A1(n5114), .A2(mgmtsoc_bus_errors_status[31]), .ZN(n5115) );
  oai22d1 U5470 ( .A1(n5116), .A2(n5204), .B1(n5217), .B2(n5115), .ZN(n3358)
         );
  ah01d1 U5471 ( .A(n5117), .B(mgmtsoc_bus_errors_status[30]), .CO(n5114), .S(
        n5118) );
  inv0d0 U5472 ( .I(n5118), .ZN(n5119) );
  oai22d1 U5473 ( .A1(n5120), .A2(n5204), .B1(n5217), .B2(n5119), .ZN(n3357)
         );
  buffd1 U5474 ( .I(n5204), .Z(n5238) );
  ah01d1 U5475 ( .A(n5121), .B(mgmtsoc_bus_errors_status[29]), .CO(n5117), .S(
        n5122) );
  inv0d0 U5476 ( .I(n5122), .ZN(n5123) );
  oai22d1 U5477 ( .A1(n5124), .A2(n5238), .B1(n5217), .B2(n5123), .ZN(n3356)
         );
  ah01d1 U5478 ( .A(n5125), .B(mgmtsoc_bus_errors_status[28]), .CO(n5121), .S(
        n5126) );
  inv0d0 U5479 ( .I(n5126), .ZN(n5127) );
  oai22d1 U5480 ( .A1(n5128), .A2(n5238), .B1(n5217), .B2(n5127), .ZN(n3355)
         );
  ah01d1 U5481 ( .A(n5129), .B(mgmtsoc_bus_errors_status[27]), .CO(n5125), .S(
        n5130) );
  inv0d0 U5482 ( .I(n5130), .ZN(n5131) );
  oai22d1 U5483 ( .A1(n5132), .A2(n5204), .B1(n5217), .B2(n5131), .ZN(n3354)
         );
  ah01d1 U5484 ( .A(n5133), .B(mgmtsoc_bus_errors_status[26]), .CO(n5129), .S(
        n5134) );
  inv0d0 U5485 ( .I(n5134), .ZN(n5135) );
  oai22d1 U5486 ( .A1(n5136), .A2(n5204), .B1(n5217), .B2(n5135), .ZN(n3353)
         );
  ah01d1 U5487 ( .A(n5137), .B(mgmtsoc_bus_errors_status[25]), .CO(n5133), .S(
        n5138) );
  inv0d0 U5488 ( .I(n5138), .ZN(n5139) );
  oai22d1 U5489 ( .A1(n5140), .A2(n5204), .B1(n5217), .B2(n5139), .ZN(n3352)
         );
  ah01d1 U5490 ( .A(n5141), .B(mgmtsoc_bus_errors_status[24]), .CO(n5137), .S(
        n5142) );
  inv0d0 U5491 ( .I(n5142), .ZN(n5143) );
  oai22d1 U5492 ( .A1(n5144), .A2(n5238), .B1(n5217), .B2(n5143), .ZN(n3351)
         );
  buffd1 U5493 ( .I(n5217), .Z(n5237) );
  ah01d1 U5494 ( .A(n5145), .B(mgmtsoc_bus_errors_status[23]), .CO(n5141), .S(
        n5146) );
  inv0d0 U5495 ( .I(n5146), .ZN(n5147) );
  oai22d1 U5496 ( .A1(n5148), .A2(n5204), .B1(n5237), .B2(n5147), .ZN(n3350)
         );
  ah01d1 U5497 ( .A(n5149), .B(mgmtsoc_bus_errors_status[22]), .CO(n5145), .S(
        n5150) );
  inv0d0 U5498 ( .I(n5150), .ZN(n5151) );
  oai22d1 U5499 ( .A1(n5152), .A2(n5238), .B1(n5217), .B2(n5151), .ZN(n3349)
         );
  ah01d1 U5500 ( .A(n5153), .B(mgmtsoc_bus_errors_status[21]), .CO(n5149), .S(
        n5154) );
  inv0d0 U5501 ( .I(n5154), .ZN(n5155) );
  oai22d1 U5502 ( .A1(n5156), .A2(n5238), .B1(n5217), .B2(n5155), .ZN(n3348)
         );
  ah01d1 U5503 ( .A(n5157), .B(mgmtsoc_bus_errors_status[20]), .CO(n5153), .S(
        n5158) );
  inv0d0 U5504 ( .I(n5158), .ZN(n5159) );
  oai22d1 U5505 ( .A1(n5160), .A2(n5204), .B1(n5237), .B2(n5159), .ZN(n3347)
         );
  ah01d1 U5506 ( .A(n5161), .B(mgmtsoc_bus_errors_status[19]), .CO(n5157), .S(
        n5162) );
  inv0d0 U5507 ( .I(n5162), .ZN(n5163) );
  oai22d1 U5508 ( .A1(n5164), .A2(n5238), .B1(n5217), .B2(n5163), .ZN(n3346)
         );
  ah01d1 U5509 ( .A(n5165), .B(mgmtsoc_bus_errors_status[18]), .CO(n5161), .S(
        n5166) );
  inv0d0 U5510 ( .I(n5166), .ZN(n5167) );
  oai22d1 U5511 ( .A1(n5168), .A2(n5204), .B1(n5237), .B2(n5167), .ZN(n3345)
         );
  ah01d1 U5512 ( .A(n5169), .B(mgmtsoc_bus_errors_status[17]), .CO(n5165), .S(
        n5170) );
  inv0d0 U5513 ( .I(n5170), .ZN(n5171) );
  oai22d1 U5514 ( .A1(n5172), .A2(n5238), .B1(n5237), .B2(n5171), .ZN(n3344)
         );
  ah01d1 U5515 ( .A(n5173), .B(mgmtsoc_bus_errors_status[16]), .CO(n5169), .S(
        n5174) );
  inv0d0 U5516 ( .I(n5174), .ZN(n5175) );
  oai22d1 U5517 ( .A1(n5176), .A2(n5204), .B1(n5237), .B2(n5175), .ZN(n3343)
         );
  ah01d1 U5518 ( .A(n5177), .B(mgmtsoc_bus_errors_status[15]), .CO(n5173), .S(
        n5178) );
  inv0d0 U5519 ( .I(n5178), .ZN(n5179) );
  oai22d1 U5520 ( .A1(n5180), .A2(n5238), .B1(n5237), .B2(n5179), .ZN(n3342)
         );
  ah01d1 U5521 ( .A(n5181), .B(mgmtsoc_bus_errors_status[14]), .CO(n5177), .S(
        n5182) );
  inv0d0 U5522 ( .I(n5182), .ZN(n5183) );
  oai22d1 U5523 ( .A1(n5184), .A2(n5204), .B1(n5237), .B2(n5183), .ZN(n3341)
         );
  ah01d1 U5524 ( .A(n5185), .B(mgmtsoc_bus_errors_status[13]), .CO(n5181), .S(
        n5186) );
  inv0d0 U5525 ( .I(n5186), .ZN(n5187) );
  oai22d1 U5526 ( .A1(n5188), .A2(n5204), .B1(n5237), .B2(n5187), .ZN(n3340)
         );
  ah01d1 U5527 ( .A(n5189), .B(mgmtsoc_bus_errors_status[12]), .CO(n5185), .S(
        n5190) );
  inv0d0 U5528 ( .I(n5190), .ZN(n5191) );
  oai22d1 U5529 ( .A1(n5192), .A2(n5204), .B1(n5237), .B2(n5191), .ZN(n3339)
         );
  ah01d1 U5530 ( .A(n5193), .B(mgmtsoc_bus_errors_status[11]), .CO(n5189), .S(
        n5194) );
  inv0d0 U5531 ( .I(n5194), .ZN(n5195) );
  oai22d1 U5532 ( .A1(n5196), .A2(n5204), .B1(n5237), .B2(n5195), .ZN(n3338)
         );
  ah01d1 U5533 ( .A(n5197), .B(mgmtsoc_bus_errors_status[10]), .CO(n5193), .S(
        n5198) );
  inv0d0 U5534 ( .I(n5198), .ZN(n5199) );
  oai22d1 U5535 ( .A1(n5200), .A2(n5238), .B1(n5217), .B2(n5199), .ZN(n3337)
         );
  ah01d1 U5536 ( .A(n5201), .B(mgmtsoc_bus_errors_status[9]), .CO(n5197), .S(
        n5202) );
  inv0d0 U5537 ( .I(n5202), .ZN(n5203) );
  oai22d1 U5538 ( .A1(n5205), .A2(n5204), .B1(n5237), .B2(n5203), .ZN(n3336)
         );
  ah01d1 U5539 ( .A(n5206), .B(mgmtsoc_bus_errors_status[8]), .CO(n5201), .S(
        n5207) );
  inv0d0 U5540 ( .I(n5207), .ZN(n5208) );
  oai22d1 U5541 ( .A1(n5209), .A2(n5238), .B1(n5217), .B2(n5208), .ZN(n3335)
         );
  ah01d1 U5542 ( .A(n5210), .B(mgmtsoc_bus_errors_status[7]), .CO(n5206), .S(
        n5211) );
  inv0d0 U5543 ( .I(n5211), .ZN(n5212) );
  oai22d1 U5544 ( .A1(n5213), .A2(n5238), .B1(n5237), .B2(n5212), .ZN(n3334)
         );
  ah01d1 U5545 ( .A(n5214), .B(mgmtsoc_bus_errors_status[6]), .CO(n5210), .S(
        n5215) );
  inv0d0 U5546 ( .I(n5215), .ZN(n5216) );
  oai22d1 U5547 ( .A1(n5218), .A2(n5238), .B1(n5217), .B2(n5216), .ZN(n3333)
         );
  ah01d1 U5548 ( .A(n5219), .B(mgmtsoc_bus_errors_status[5]), .CO(n5214), .S(
        n5220) );
  inv0d0 U5549 ( .I(n5220), .ZN(n5221) );
  oai22d1 U5550 ( .A1(n5222), .A2(n5238), .B1(n5237), .B2(n5221), .ZN(n3332)
         );
  ah01d1 U5551 ( .A(n5223), .B(mgmtsoc_bus_errors_status[4]), .CO(n5219), .S(
        n5224) );
  inv0d0 U5552 ( .I(n5224), .ZN(n5225) );
  oai22d1 U5553 ( .A1(n5226), .A2(n5238), .B1(n5237), .B2(n5225), .ZN(n3331)
         );
  ah01d1 U5554 ( .A(n5227), .B(mgmtsoc_bus_errors_status[3]), .CO(n5223), .S(
        n5228) );
  inv0d0 U5555 ( .I(n5228), .ZN(n5229) );
  oai22d1 U5556 ( .A1(n5230), .A2(n5238), .B1(n5237), .B2(n5229), .ZN(n3330)
         );
  ah01d1 U5557 ( .A(n5231), .B(mgmtsoc_bus_errors_status[2]), .CO(n5227), .S(
        n5232) );
  inv0d0 U5558 ( .I(n5232), .ZN(n5233) );
  oai22d1 U5559 ( .A1(n5234), .A2(n5238), .B1(n5237), .B2(n5233), .ZN(n3329)
         );
  ah01d1 U5560 ( .A(mgmtsoc_bus_errors_status[0]), .B(
        mgmtsoc_bus_errors_status[1]), .CO(n5231), .S(n5235) );
  inv0d0 U5561 ( .I(n5235), .ZN(n5236) );
  oai22d1 U5562 ( .A1(n5239), .A2(n5238), .B1(n5237), .B2(n5236), .ZN(n3328)
         );
  buffd1 U5563 ( .I(n5286), .Z(n5282) );
  oaim21d1 U5564 ( .B1(n5241), .B2(n5240), .A(n4881), .ZN(n5285) );
  oai22d1 U5565 ( .A1(n4808), .A2(n5282), .B1(n5242), .B2(n5285), .ZN(n3327)
         );
  oai22d1 U5566 ( .A1(n5294), .A2(n5282), .B1(n5243), .B2(n5285), .ZN(n3326)
         );
  buffd1 U5567 ( .I(n5285), .Z(n5279) );
  oai22d1 U5568 ( .A1(n5245), .A2(n5282), .B1(n5279), .B2(n5244), .ZN(n3325)
         );
  inv0d1 U5569 ( .I(n5282), .ZN(n5277) );
  aoim22d1 U5570 ( .A1(n5277), .A2(n5246), .B1(csrbank0_scratch0_w[3]), .B2(
        n5279), .Z(n3324) );
  aoim22d1 U5571 ( .A1(n5277), .A2(n5247), .B1(csrbank0_scratch0_w[4]), .B2(
        n5279), .Z(n3323) );
  aoim22d1 U5572 ( .A1(n5277), .A2(n5248), .B1(csrbank0_scratch0_w[5]), .B2(
        n5285), .Z(n3322) );
  aoim22d1 U5573 ( .A1(n5277), .A2(n5249), .B1(csrbank0_scratch0_w[6]), .B2(
        n5279), .Z(n3321) );
  oai22d1 U5574 ( .A1(n5251), .A2(n5282), .B1(n5285), .B2(n5250), .ZN(n3320)
         );
  oai22d1 U5575 ( .A1(n4783), .A2(n5282), .B1(n5285), .B2(n5252), .ZN(n3319)
         );
  aoim22d1 U5576 ( .A1(n5277), .A2(n4593), .B1(csrbank0_scratch0_w[9]), .B2(
        n5279), .Z(n3318) );
  aoim22d1 U5577 ( .A1(n5277), .A2(n4595), .B1(csrbank0_scratch0_w[10]), .B2(
        n5279), .Z(n3317) );
  oai22d1 U5578 ( .A1(n5254), .A2(n5282), .B1(n5279), .B2(n5253), .ZN(n3316)
         );
  aoim22d1 U5579 ( .A1(n5277), .A2(n4598), .B1(csrbank0_scratch0_w[12]), .B2(
        n5285), .Z(n3315) );
  oai22d1 U5580 ( .A1(n4790), .A2(n5286), .B1(n5285), .B2(n5255), .ZN(n3314)
         );
  aoim22d1 U5581 ( .A1(n5277), .A2(n4601), .B1(csrbank0_scratch0_w[14]), .B2(
        n5279), .Z(n3313) );
  oai22d1 U5582 ( .A1(n4793), .A2(n5286), .B1(n5285), .B2(n5256), .ZN(n3312)
         );
  oai22d1 U5583 ( .A1(n2003), .A2(n5286), .B1(n5279), .B2(n5257), .ZN(n3311)
         );
  oai22d1 U5584 ( .A1(n5259), .A2(n5282), .B1(n5279), .B2(n5258), .ZN(n3310)
         );
  aoim22d1 U5585 ( .A1(n5277), .A2(n5260), .B1(csrbank0_scratch0_w[18]), .B2(
        n5285), .Z(n3309) );
  oai22d1 U5586 ( .A1(n5262), .A2(n5282), .B1(n5285), .B2(n5261), .ZN(n3308)
         );
  aoim22d1 U5587 ( .A1(n5277), .A2(n5263), .B1(csrbank0_scratch0_w[20]), .B2(
        n5285), .Z(n3307) );
  aoim22d1 U5588 ( .A1(n5277), .A2(n5264), .B1(csrbank0_scratch0_w[21]), .B2(
        n5285), .Z(n3306) );
  oai22d1 U5589 ( .A1(n5266), .A2(n5286), .B1(n5285), .B2(n5265), .ZN(n3305)
         );
  oai22d1 U5590 ( .A1(n5268), .A2(n5282), .B1(n5279), .B2(n5267), .ZN(n3304)
         );
  oai22d1 U5591 ( .A1(n5270), .A2(n5286), .B1(n5285), .B2(n5269), .ZN(n3303)
         );
  aoim22d1 U5592 ( .A1(n5277), .A2(n5271), .B1(csrbank0_scratch0_w[25]), .B2(
        n5279), .Z(n3302) );
  oai22d1 U5593 ( .A1(n5273), .A2(n5282), .B1(n5279), .B2(n5272), .ZN(n3301)
         );
  oai22d1 U5594 ( .A1(n5275), .A2(n5286), .B1(n5279), .B2(n5274), .ZN(n3300)
         );
  aoim22d1 U5595 ( .A1(n5277), .A2(n5276), .B1(csrbank0_scratch0_w[28]), .B2(
        n5279), .Z(n3299) );
  oai22d1 U5596 ( .A1(n5280), .A2(n5286), .B1(n5279), .B2(n5278), .ZN(n3298)
         );
  oai22d1 U5597 ( .A1(n5283), .A2(n5282), .B1(n5285), .B2(n5281), .ZN(n3297)
         );
  oai22d1 U5598 ( .A1(n5287), .A2(n5286), .B1(n5285), .B2(n5284), .ZN(n3296)
         );
  inv0d0 U5599 ( .I(N5168), .ZN(n5293) );
  nd02d0 U5600 ( .A1(n5288), .A2(n5293), .ZN(n5291) );
  oai22d1 U5601 ( .A1(n5290), .A2(n5293), .B1(n5289), .B2(n5291), .ZN(n3295)
         );
  oai22d1 U5602 ( .A1(n5294), .A2(n5293), .B1(n5292), .B2(n5291), .ZN(n3294)
         );
  inv0d0 U5603 ( .I(n5318), .ZN(n5295) );
  aoi31d1 U5604 ( .B1(n5297), .B2(n5488), .B3(n5296), .A(n5295), .ZN(n5298) );
  oai21d1 U5605 ( .B1(n5300), .B2(n5299), .A(n5298), .ZN(n5302) );
  an02d0 U5606 ( .A1(n5340), .A2(n5491), .Z(n5592) );
  buffd1 U5607 ( .I(n5592), .Z(n5604) );
  aoim22d1 U5608 ( .A1(dbg_uart_words_count[0]), .A2(n5302), .B1(n5604), .B2(
        dbg_uart_words_count[0]), .Z(n3293) );
  inv0d0 U5609 ( .I(n5302), .ZN(n5315) );
  aor22d1 U5610 ( .A1(n5604), .A2(n5303), .B1(n5315), .B2(
        dbg_uart_words_count[1]), .Z(n3292) );
  ah01d1 U5611 ( .A(dbg_uart_words_count[0]), .B(dbg_uart_words_count[1]), 
        .CO(n5305), .S(n5303) );
  aor22d1 U5612 ( .A1(n5604), .A2(n5304), .B1(n5315), .B2(
        dbg_uart_words_count[2]), .Z(n3291) );
  ah01d1 U5613 ( .A(n5305), .B(dbg_uart_words_count[2]), .CO(n5307), .S(n5304)
         );
  aor22d1 U5614 ( .A1(n5604), .A2(n5306), .B1(n5315), .B2(
        dbg_uart_words_count[3]), .Z(n3290) );
  ah01d1 U5615 ( .A(n5307), .B(dbg_uart_words_count[3]), .CO(n5309), .S(n5306)
         );
  aor22d1 U5616 ( .A1(n5604), .A2(n5308), .B1(n5315), .B2(
        dbg_uart_words_count[4]), .Z(n3289) );
  ah01d1 U5617 ( .A(n5309), .B(dbg_uart_words_count[4]), .CO(n5311), .S(n5308)
         );
  aor22d1 U5618 ( .A1(n5604), .A2(n5310), .B1(n5315), .B2(
        dbg_uart_words_count[5]), .Z(n3288) );
  ah01d1 U5619 ( .A(n5311), .B(dbg_uart_words_count[5]), .CO(n5313), .S(n5310)
         );
  aor22d1 U5620 ( .A1(n5604), .A2(n5312), .B1(n5315), .B2(
        dbg_uart_words_count[6]), .Z(n3287) );
  ah01d1 U5621 ( .A(n5313), .B(dbg_uart_words_count[6]), .CO(n5314), .S(n5312)
         );
  xr02d1 U5622 ( .A1(n5314), .A2(dbg_uart_words_count[7]), .Z(n5316) );
  aor22d1 U5623 ( .A1(n5604), .A2(n5316), .B1(n5315), .B2(
        dbg_uart_words_count[7]), .Z(n3286) );
  inv0d0 U5624 ( .I(n5342), .ZN(n5326) );
  nr02d0 U5625 ( .A1(n5326), .A2(n5320), .ZN(n5317) );
  nd02d0 U5626 ( .A1(n5318), .A2(n5317), .ZN(n5322) );
  oai21d1 U5627 ( .B1(n5326), .B2(n5320), .A(n5319), .ZN(n5324) );
  inv0d0 U5628 ( .I(dbg_uart_bytes_count[0]), .ZN(n5321) );
  aoi22d1 U5629 ( .A1(dbg_uart_bytes_count[0]), .A2(n5322), .B1(n5324), .B2(
        n5321), .ZN(n3285) );
  nr02d0 U5630 ( .A1(dbg_uart_bytes_count[1]), .A2(n5321), .ZN(n6012) );
  inv0d0 U5631 ( .I(dbg_uart_bytes_count[1]), .ZN(n5323) );
  nr02d0 U5632 ( .A1(dbg_uart_bytes_count[0]), .A2(n5323), .ZN(n6013) );
  nr02d0 U5633 ( .A1(n6012), .A2(n6013), .ZN(n5325) );
  oai22d1 U5634 ( .A1(n5325), .A2(n5324), .B1(n5323), .B2(n5322), .ZN(n3284)
         );
  nd03d1 U5635 ( .A1(uartwishbonebridge_state[0]), .A2(n5326), .A3(n5956), 
        .ZN(n5482) );
  nr02d0 U5636 ( .A1(n5341), .A2(n5488), .ZN(n5327) );
  nr04d0 U5637 ( .A1(interface9_bank_bus_dat_r[0]), .A2(
        \interface7_bank_bus_dat_r[0] ), .A3(\interface14_bank_bus_dat_r[0] ), 
        .A4(interface11_bank_bus_dat_r[0]), .ZN(n5338) );
  nr04d0 U5638 ( .A1(\interface2_bank_bus_dat_r[0] ), .A2(
        \interface12_bank_bus_dat_r[0] ), .A3(\interface13_bank_bus_dat_r[0] ), 
        .A4(interface19_bank_bus_dat_r[0]), .ZN(n5331) );
  nr04d0 U5639 ( .A1(\interface15_bank_bus_dat_r[0] ), .A2(
        \interface16_bank_bus_dat_r[0] ), .A3(\interface17_bank_bus_dat_r[0] ), 
        .A4(\interface18_bank_bus_dat_r[0] ), .ZN(n5330) );
  nr04d0 U5640 ( .A1(interface10_bank_bus_dat_r[0]), .A2(
        interface0_bank_bus_dat_r[0]), .A3(\interface5_bank_bus_dat_r[0] ), 
        .A4(interface6_bank_bus_dat_r[0]), .ZN(n5329) );
  nr04d0 U5641 ( .A1(interface3_bank_bus_dat_r[0]), .A2(
        \interface1_bank_bus_dat_r[0] ), .A3(\interface8_bank_bus_dat_r[0] ), 
        .A4(interface4_bank_bus_dat_r[0]), .ZN(n5328) );
  an04d0 U5642 ( .A1(n5331), .A2(n5330), .A3(n5329), .A4(n5328), .Z(n5337) );
  aoi22d1 U5643 ( .A1(n5394), .A2(mprj_dat_i[0]), .B1(n5395), .B2(
        mgmtsoc_vexriscv_debug_bus_dat_r[0]), .ZN(n5333) );
  aoi22d1 U5644 ( .A1(n5429), .A2(hk_dat_i[0]), .B1(n5406), .B2(
        dff2_bus_dat_r[0]), .ZN(n5332) );
  oai211d1 U5645 ( .C1(n5763), .C2(n5432), .A(n5333), .B(n5332), .ZN(n5334) );
  aoi211d1 U5646 ( .C1(n1409), .C2(\RAM256/Do0_pre[0][0] ), .A(n5335), .B(
        n5334), .ZN(n5336) );
  aon211d1 U5647 ( .C1(n5338), .C2(n5337), .B(n5356), .A(n5336), .ZN(n5339) );
  aoi31d1 U5648 ( .B1(slave_sel_r[1]), .B2(\RAM256/Do0_pre[1][0] ), .B3(
        mprj_adr_o[9]), .A(n5339), .ZN(n5343) );
  inv0d0 U5649 ( .I(dbg_uart_wishbone_dat_w[0]), .ZN(n5381) );
  aon211d1 U5650 ( .C1(n5342), .C2(n5341), .B(n5488), .A(n4881), .ZN(n5487) );
  buffd1 U5651 ( .I(n5487), .Z(n5481) );
  oai222d1 U5652 ( .A1(n5482), .A2(n5969), .B1(n5467), .B2(n5343), .C1(n5381), 
        .C2(n5481), .ZN(n3283) );
  inv0d0 U5653 ( .I(n5343), .ZN(mgmtsoc_ibus_ibus_dat_r[0]) );
  buffd1 U5654 ( .I(n5482), .Z(n5452) );
  inv0d0 U5655 ( .I(mgmtsoc_ibus_ibus_dat_r[1]), .ZN(n5344) );
  inv0d0 U5656 ( .I(dbg_uart_wishbone_dat_w[1]), .ZN(n5390) );
  oai222d1 U5657 ( .A1(n5970), .A2(n5452), .B1(n5467), .B2(n5344), .C1(n5390), 
        .C2(n5481), .ZN(n3282) );
  inv0d0 U5658 ( .I(mgmtsoc_ibus_ibus_dat_r[2]), .ZN(n5345) );
  inv0d0 U5659 ( .I(dbg_uart_wishbone_dat_w[2]), .ZN(n5402) );
  oai222d1 U5660 ( .A1(n5971), .A2(n5452), .B1(n5467), .B2(n5345), .C1(n5402), 
        .C2(n5481), .ZN(n3281) );
  nr04d0 U5661 ( .A1(interface9_bank_bus_dat_r[3]), .A2(
        interface10_bank_bus_dat_r[3]), .A3(interface0_bank_bus_dat_r[3]), 
        .A4(interface11_bank_bus_dat_r[3]), .ZN(n5347) );
  aon211d1 U5662 ( .C1(n5347), .C2(n5346), .B(n5356), .A(n5425), .ZN(n5351) );
  aoi22d1 U5663 ( .A1(slave_sel_r[0]), .A2(mgmtsoc_vexriscv_debug_bus_dat_r[3]), .B1(n5429), .B2(hk_dat_i[3]), .ZN(n5349) );
  aoi22d1 U5664 ( .A1(n5394), .A2(mprj_dat_i[3]), .B1(n5406), .B2(
        dff2_bus_dat_r[3]), .ZN(n5348) );
  oai211d1 U5665 ( .C1(n5769), .C2(n5432), .A(n5349), .B(n5348), .ZN(n5350) );
  aoi211d1 U5666 ( .C1(n5435), .C2(\RAM256/Do0_pre[0][3] ), .A(n5351), .B(
        n5350), .ZN(n5352) );
  oaim21d1 U5667 ( .B1(n5437), .B2(\RAM256/Do0_pre[1][3] ), .A(n5352), .ZN(
        mgmtsoc_ibus_ibus_dat_r[3]) );
  inv0d0 U5668 ( .I(mgmtsoc_ibus_ibus_dat_r[3]), .ZN(n5353) );
  inv0d0 U5669 ( .I(dbg_uart_wishbone_dat_w[3]), .ZN(n5412) );
  oai222d1 U5670 ( .A1(n5972), .A2(n5452), .B1(n5467), .B2(n5353), .C1(n5412), 
        .C2(n5481), .ZN(n3280) );
  inv0d0 U5671 ( .I(mgmtsoc_ibus_ibus_dat_r[4]), .ZN(n5354) );
  inv0d0 U5672 ( .I(dbg_uart_wishbone_dat_w[4]), .ZN(n5414) );
  oai222d1 U5673 ( .A1(n5973), .A2(n5482), .B1(n5467), .B2(n5354), .C1(n5414), 
        .C2(n5481), .ZN(n3279) );
  buffd1 U5674 ( .I(n5467), .Z(n5485) );
  inv0d0 U5675 ( .I(mgmtsoc_ibus_ibus_dat_r[5]), .ZN(n5355) );
  inv0d0 U5676 ( .I(dbg_uart_wishbone_dat_w[5]), .ZN(n5423) );
  oai222d1 U5677 ( .A1(n5974), .A2(n5452), .B1(n5485), .B2(n5355), .C1(n5423), 
        .C2(n5487), .ZN(n3278) );
  nr04d0 U5678 ( .A1(interface9_bank_bus_dat_r[6]), .A2(
        interface10_bank_bus_dat_r[6]), .A3(interface0_bank_bus_dat_r[6]), 
        .A4(interface11_bank_bus_dat_r[6]), .ZN(n5358) );
  nr03d0 U5679 ( .A1(interface3_bank_bus_dat_r[6]), .A2(
        interface6_bank_bus_dat_r[6]), .A3(interface4_bank_bus_dat_r[6]), .ZN(
        n5357) );
  aon211d1 U5680 ( .C1(n5358), .C2(n5357), .B(n5356), .A(n5425), .ZN(n5362) );
  aoi22d1 U5681 ( .A1(n5394), .A2(mprj_dat_i[6]), .B1(n5406), .B2(
        dff2_bus_dat_r[6]), .ZN(n5360) );
  aoi22d1 U5682 ( .A1(n5395), .A2(mgmtsoc_vexriscv_debug_bus_dat_r[6]), .B1(
        n5429), .B2(hk_dat_i[6]), .ZN(n5359) );
  oai211d1 U5683 ( .C1(n5771), .C2(n5432), .A(n5360), .B(n5359), .ZN(n5361) );
  aoi211d1 U5684 ( .C1(n5437), .C2(\RAM256/Do0_pre[1][6] ), .A(n5362), .B(
        n5361), .ZN(n5363) );
  oaim21d1 U5685 ( .B1(n1409), .B2(\RAM256/Do0_pre[0][6] ), .A(n5363), .ZN(
        mgmtsoc_ibus_ibus_dat_r[6]) );
  inv0d0 U5686 ( .I(mgmtsoc_ibus_ibus_dat_r[6]), .ZN(n5364) );
  inv0d0 U5687 ( .I(dbg_uart_wishbone_dat_w[6]), .ZN(n5438) );
  oai222d1 U5688 ( .A1(n5975), .A2(n5452), .B1(n5467), .B2(n5364), .C1(n5438), 
        .C2(n5481), .ZN(n3277) );
  nr04d0 U5689 ( .A1(interface9_bank_bus_dat_r[7]), .A2(
        interface10_bank_bus_dat_r[7]), .A3(interface0_bank_bus_dat_r[7]), 
        .A4(interface11_bank_bus_dat_r[7]), .ZN(n5366) );
  aon211d1 U5690 ( .C1(n5366), .C2(n5365), .B(n5426), .A(n5425), .ZN(n5370) );
  aoi22d1 U5691 ( .A1(n5394), .A2(mprj_dat_i[7]), .B1(slave_sel_r[0]), .B2(
        mgmtsoc_vexriscv_debug_bus_dat_r[7]), .ZN(n5368) );
  aoi22d1 U5692 ( .A1(n5429), .A2(hk_dat_i[7]), .B1(n5406), .B2(
        dff2_bus_dat_r[7]), .ZN(n5367) );
  oai211d1 U5693 ( .C1(n5775), .C2(n5432), .A(n5368), .B(n5367), .ZN(n5369) );
  aoi211d1 U5694 ( .C1(n5437), .C2(\RAM256/Do0_pre[1][7] ), .A(n5370), .B(
        n5369), .ZN(n5371) );
  oaim21d1 U5695 ( .B1(n1409), .B2(\RAM256/Do0_pre[0][7] ), .A(n5371), .ZN(
        mgmtsoc_ibus_ibus_dat_r[7]) );
  inv0d0 U5696 ( .I(mgmtsoc_ibus_ibus_dat_r[7]), .ZN(n5372) );
  inv0d0 U5697 ( .I(dbg_uart_wishbone_dat_w[7]), .ZN(n5440) );
  oai222d1 U5698 ( .A1(n5976), .A2(n5452), .B1(n5485), .B2(n5372), .C1(n5440), 
        .C2(n5487), .ZN(n3276) );
  nr04d0 U5699 ( .A1(interface6_bank_bus_dat_r[8]), .A2(
        interface3_bank_bus_dat_r[8]), .A3(interface10_bank_bus_dat_r[8]), 
        .A4(interface9_bank_bus_dat_r[8]), .ZN(n5374) );
  inv0d0 U5700 ( .I(interface0_bank_bus_dat_r[8]), .ZN(n5373) );
  aon211d1 U5701 ( .C1(n5374), .C2(n5373), .B(n5426), .A(n5425), .ZN(n5378) );
  aoi22d1 U5702 ( .A1(n5394), .A2(mprj_dat_i[8]), .B1(n5406), .B2(
        dff2_bus_dat_r[8]), .ZN(n5376) );
  aoi22d1 U5703 ( .A1(slave_sel_r[0]), .A2(mgmtsoc_vexriscv_debug_bus_dat_r[8]), .B1(slave_sel_r[5]), .B2(hk_dat_i[8]), .ZN(n5375) );
  oai211d1 U5704 ( .C1(n5755), .C2(n5432), .A(n5376), .B(n5375), .ZN(n5377) );
  aoi211d1 U5705 ( .C1(n1409), .C2(\RAM256/Do0_pre[0][8] ), .A(n5378), .B(
        n5377), .ZN(n5379) );
  oaim21d1 U5706 ( .B1(n5380), .B2(\RAM256/Do0_pre[1][8] ), .A(n5379), .ZN(
        mgmtsoc_ibus_ibus_dat_r[8]) );
  inv0d0 U5707 ( .I(dbg_uart_wishbone_dat_w[8]), .ZN(n5442) );
  inv0d0 U5708 ( .I(mgmtsoc_ibus_ibus_dat_r[8]), .ZN(n5382) );
  oai222d1 U5709 ( .A1(n5487), .A2(n5442), .B1(n5467), .B2(n5382), .C1(n5381), 
        .C2(n5452), .ZN(n3275) );
  nr04d0 U5710 ( .A1(interface6_bank_bus_dat_r[9]), .A2(
        interface3_bank_bus_dat_r[9]), .A3(interface10_bank_bus_dat_r[9]), 
        .A4(interface9_bank_bus_dat_r[9]), .ZN(n5384) );
  inv0d0 U5711 ( .I(interface0_bank_bus_dat_r[9]), .ZN(n5383) );
  aon211d1 U5712 ( .C1(n5384), .C2(n5383), .B(n5426), .A(n5425), .ZN(n5388) );
  aoi22d1 U5713 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[9]), .B1(slave_sel_r[2]), 
        .B2(dff2_bus_dat_r[9]), .ZN(n5386) );
  aoi22d1 U5714 ( .A1(n5395), .A2(mgmtsoc_vexriscv_debug_bus_dat_r[9]), .B1(
        slave_sel_r[5]), .B2(hk_dat_i[9]), .ZN(n5385) );
  oai211d1 U5715 ( .C1(n5756), .C2(n5432), .A(n5386), .B(n5385), .ZN(n5387) );
  aoi211d1 U5716 ( .C1(n5437), .C2(\RAM256/Do0_pre[1][9] ), .A(n5388), .B(
        n5387), .ZN(n5389) );
  oaim21d1 U5717 ( .B1(n1409), .B2(\RAM256/Do0_pre[0][9] ), .A(n5389), .ZN(
        mgmtsoc_ibus_ibus_dat_r[9]) );
  inv0d0 U5718 ( .I(dbg_uart_wishbone_dat_w[9]), .ZN(n5444) );
  inv0d0 U5719 ( .I(mgmtsoc_ibus_ibus_dat_r[9]), .ZN(n5391) );
  oai222d1 U5720 ( .A1(n5481), .A2(n5444), .B1(n5485), .B2(n5391), .C1(n5390), 
        .C2(n5452), .ZN(n3274) );
  inv0d0 U5721 ( .I(interface0_bank_bus_dat_r[10]), .ZN(n5392) );
  aon211d1 U5722 ( .C1(n5393), .C2(n5392), .B(n5426), .A(n5425), .ZN(n5399) );
  aoi22d1 U5723 ( .A1(n5394), .A2(mprj_dat_i[10]), .B1(n5406), .B2(
        dff2_bus_dat_r[10]), .ZN(n5397) );
  aoi22d1 U5724 ( .A1(n5395), .A2(mgmtsoc_vexriscv_debug_bus_dat_r[10]), .B1(
        slave_sel_r[5]), .B2(hk_dat_i[10]), .ZN(n5396) );
  oai211d1 U5725 ( .C1(n5757), .C2(n5432), .A(n5397), .B(n5396), .ZN(n5398) );
  aoi211d1 U5726 ( .C1(n5435), .C2(\RAM256/Do0_pre[0][10] ), .A(n5399), .B(
        n5398), .ZN(n5400) );
  oaim21d1 U5727 ( .B1(n5401), .B2(\RAM256/Do0_pre[1][10] ), .A(n5400), .ZN(
        mgmtsoc_ibus_ibus_dat_r[10]) );
  inv0d0 U5728 ( .I(dbg_uart_wishbone_dat_w[10]), .ZN(n5446) );
  inv0d0 U5729 ( .I(mgmtsoc_ibus_ibus_dat_r[10]), .ZN(n5403) );
  oai222d1 U5730 ( .A1(n5487), .A2(n5446), .B1(n5467), .B2(n5403), .C1(n5402), 
        .C2(n5452), .ZN(n3273) );
  nr04d0 U5731 ( .A1(interface6_bank_bus_dat_r[11]), .A2(
        interface3_bank_bus_dat_r[11]), .A3(interface10_bank_bus_dat_r[11]), 
        .A4(interface9_bank_bus_dat_r[11]), .ZN(n5405) );
  inv0d0 U5732 ( .I(interface0_bank_bus_dat_r[11]), .ZN(n5404) );
  aon211d1 U5733 ( .C1(n5405), .C2(n5404), .B(n5426), .A(n5425), .ZN(n5410) );
  aoi22d1 U5734 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[11]), .B1(n5406), .B2(
        dff2_bus_dat_r[11]), .ZN(n5408) );
  aoi22d1 U5735 ( .A1(slave_sel_r[0]), .A2(
        mgmtsoc_vexriscv_debug_bus_dat_r[11]), .B1(slave_sel_r[5]), .B2(
        hk_dat_i[11]), .ZN(n5407) );
  oai211d1 U5736 ( .C1(n5758), .C2(n5432), .A(n5408), .B(n5407), .ZN(n5409) );
  aoi211d1 U5737 ( .C1(n5435), .C2(\RAM256/Do0_pre[0][11] ), .A(n5410), .B(
        n5409), .ZN(n5411) );
  oaim21d1 U5738 ( .B1(n5437), .B2(\RAM256/Do0_pre[1][11] ), .A(n5411), .ZN(
        mgmtsoc_ibus_ibus_dat_r[11]) );
  inv0d0 U5739 ( .I(dbg_uart_wishbone_dat_w[11]), .ZN(n5448) );
  inv0d0 U5740 ( .I(mgmtsoc_ibus_ibus_dat_r[11]), .ZN(n5413) );
  oai222d1 U5741 ( .A1(n5487), .A2(n5448), .B1(n5485), .B2(n5413), .C1(n5412), 
        .C2(n5452), .ZN(n3272) );
  inv0d0 U5742 ( .I(dbg_uart_wishbone_dat_w[12]), .ZN(n5450) );
  inv0d0 U5743 ( .I(mgmtsoc_ibus_ibus_dat_r[12]), .ZN(n5415) );
  oai222d1 U5744 ( .A1(n5481), .A2(n5450), .B1(n5485), .B2(n5415), .C1(n5414), 
        .C2(n5452), .ZN(n3271) );
  nr04d0 U5745 ( .A1(interface6_bank_bus_dat_r[13]), .A2(
        interface3_bank_bus_dat_r[13]), .A3(interface10_bank_bus_dat_r[13]), 
        .A4(interface9_bank_bus_dat_r[13]), .ZN(n5417) );
  inv0d0 U5746 ( .I(interface0_bank_bus_dat_r[13]), .ZN(n5416) );
  aon211d1 U5747 ( .C1(n5417), .C2(n5416), .B(n5426), .A(n5425), .ZN(n5421) );
  aoi22d1 U5748 ( .A1(slave_sel_r[0]), .A2(
        mgmtsoc_vexriscv_debug_bus_dat_r[13]), .B1(slave_sel_r[5]), .B2(
        hk_dat_i[13]), .ZN(n5419) );
  aoi22d1 U5749 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[13]), .B1(slave_sel_r[2]), .B2(dff2_bus_dat_r[13]), .ZN(n5418) );
  oai211d1 U5750 ( .C1(n5760), .C2(n5432), .A(n5419), .B(n5418), .ZN(n5420) );
  aoi211d1 U5751 ( .C1(n5435), .C2(\RAM256/Do0_pre[0][13] ), .A(n5421), .B(
        n5420), .ZN(n5422) );
  oaim21d1 U5752 ( .B1(n5437), .B2(\RAM256/Do0_pre[1][13] ), .A(n5422), .ZN(
        mgmtsoc_ibus_ibus_dat_r[13]) );
  inv0d0 U5753 ( .I(dbg_uart_wishbone_dat_w[13]), .ZN(n5453) );
  inv0d0 U5754 ( .I(mgmtsoc_ibus_ibus_dat_r[13]), .ZN(n5424) );
  oai222d1 U5755 ( .A1(n5487), .A2(n5453), .B1(n5485), .B2(n5424), .C1(n5423), 
        .C2(n5452), .ZN(n3270) );
  inv0d0 U5756 ( .I(interface0_bank_bus_dat_r[14]), .ZN(n5427) );
  aon211d1 U5757 ( .C1(n5428), .C2(n5427), .B(n5426), .A(n5425), .ZN(n5434) );
  aoi22d1 U5758 ( .A1(slave_sel_r[4]), .A2(mprj_dat_i[14]), .B1(slave_sel_r[2]), .B2(dff2_bus_dat_r[14]), .ZN(n5431) );
  aoi22d1 U5759 ( .A1(slave_sel_r[0]), .A2(
        mgmtsoc_vexriscv_debug_bus_dat_r[14]), .B1(n5429), .B2(hk_dat_i[14]), 
        .ZN(n5430) );
  oai211d1 U5760 ( .C1(n5761), .C2(n5432), .A(n5431), .B(n5430), .ZN(n5433) );
  aoi211d1 U5761 ( .C1(n5435), .C2(\RAM256/Do0_pre[0][14] ), .A(n5434), .B(
        n5433), .ZN(n5436) );
  oaim21d1 U5762 ( .B1(n5437), .B2(\RAM256/Do0_pre[1][14] ), .A(n5436), .ZN(
        mgmtsoc_ibus_ibus_dat_r[14]) );
  inv0d0 U5763 ( .I(dbg_uart_wishbone_dat_w[14]), .ZN(n5455) );
  inv0d0 U5764 ( .I(mgmtsoc_ibus_ibus_dat_r[14]), .ZN(n5439) );
  oai222d1 U5765 ( .A1(n5487), .A2(n5455), .B1(n5467), .B2(n5439), .C1(n5438), 
        .C2(n5452), .ZN(n3269) );
  inv0d0 U5766 ( .I(dbg_uart_wishbone_dat_w[15]), .ZN(n5457) );
  inv0d0 U5767 ( .I(mgmtsoc_ibus_ibus_dat_r[15]), .ZN(n5441) );
  oai222d1 U5768 ( .A1(n5487), .A2(n5457), .B1(n5485), .B2(n5441), .C1(n5440), 
        .C2(n5452), .ZN(n3268) );
  inv0d0 U5769 ( .I(dbg_uart_wishbone_dat_w[16]), .ZN(n5459) );
  inv0d0 U5770 ( .I(mgmtsoc_ibus_ibus_dat_r[16]), .ZN(n5443) );
  oai222d1 U5771 ( .A1(n5481), .A2(n5459), .B1(n5467), .B2(n5443), .C1(n5442), 
        .C2(n5452), .ZN(n3267) );
  inv0d0 U5772 ( .I(dbg_uart_wishbone_dat_w[17]), .ZN(n5462) );
  inv0d0 U5773 ( .I(mgmtsoc_ibus_ibus_dat_r[17]), .ZN(n5445) );
  oai222d1 U5774 ( .A1(n5487), .A2(n5462), .B1(n5485), .B2(n5445), .C1(n5444), 
        .C2(n5482), .ZN(n3266) );
  inv0d0 U5775 ( .I(dbg_uart_wishbone_dat_w[18]), .ZN(n5465) );
  inv0d0 U5776 ( .I(mgmtsoc_ibus_ibus_dat_r[18]), .ZN(n5447) );
  oai222d1 U5777 ( .A1(n5487), .A2(n5465), .B1(n5467), .B2(n5447), .C1(n5446), 
        .C2(n5452), .ZN(n3265) );
  inv0d0 U5778 ( .I(dbg_uart_wishbone_dat_w[19]), .ZN(n5469) );
  inv0d0 U5779 ( .I(mgmtsoc_ibus_ibus_dat_r[19]), .ZN(n5449) );
  oai222d1 U5780 ( .A1(n5481), .A2(n5469), .B1(n5467), .B2(n5449), .C1(n5448), 
        .C2(n5482), .ZN(n3264) );
  inv0d0 U5781 ( .I(dbg_uart_wishbone_dat_w[20]), .ZN(n5472) );
  inv0d0 U5782 ( .I(mgmtsoc_ibus_ibus_dat_r[20]), .ZN(n5451) );
  oai222d1 U5783 ( .A1(n5481), .A2(n5472), .B1(n5485), .B2(n5451), .C1(n5450), 
        .C2(n5482), .ZN(n3263) );
  inv0d0 U5784 ( .I(dbg_uart_wishbone_dat_w[21]), .ZN(n5475) );
  inv0d0 U5785 ( .I(mgmtsoc_ibus_ibus_dat_r[21]), .ZN(n5454) );
  oai222d1 U5786 ( .A1(n5487), .A2(n5475), .B1(n5485), .B2(n5454), .C1(n5453), 
        .C2(n5452), .ZN(n3262) );
  inv0d0 U5787 ( .I(dbg_uart_wishbone_dat_w[22]), .ZN(n5478) );
  inv0d0 U5788 ( .I(mgmtsoc_ibus_ibus_dat_r[22]), .ZN(n5456) );
  oai222d1 U5789 ( .A1(n5481), .A2(n5478), .B1(n5467), .B2(n5456), .C1(n5455), 
        .C2(n5482), .ZN(n3261) );
  inv0d0 U5790 ( .I(dbg_uart_wishbone_dat_w[23]), .ZN(n5483) );
  inv0d0 U5791 ( .I(mgmtsoc_ibus_ibus_dat_r[23]), .ZN(n5458) );
  oai222d1 U5792 ( .A1(n5481), .A2(n5483), .B1(n5485), .B2(n5458), .C1(n5457), 
        .C2(n5482), .ZN(n3260) );
  inv0d0 U5793 ( .I(dbg_uart_wishbone_dat_w[24]), .ZN(n5461) );
  inv0d0 U5794 ( .I(mgmtsoc_ibus_ibus_dat_r[24]), .ZN(n5460) );
  oai222d1 U5795 ( .A1(n5481), .A2(n5461), .B1(n5485), .B2(n5460), .C1(n5459), 
        .C2(n5482), .ZN(n3259) );
  inv0d0 U5796 ( .I(dbg_uart_wishbone_dat_w[25]), .ZN(n5464) );
  inv0d0 U5797 ( .I(mgmtsoc_ibus_ibus_dat_r[25]), .ZN(n5463) );
  oai222d1 U5798 ( .A1(n5481), .A2(n5464), .B1(n5467), .B2(n5463), .C1(n5462), 
        .C2(n5482), .ZN(n3258) );
  inv0d0 U5799 ( .I(dbg_uart_wishbone_dat_w[26]), .ZN(n5468) );
  inv0d0 U5800 ( .I(mgmtsoc_ibus_ibus_dat_r[26]), .ZN(n5466) );
  oai222d1 U5801 ( .A1(n5487), .A2(n5468), .B1(n5467), .B2(n5466), .C1(n5465), 
        .C2(n5482), .ZN(n3257) );
  inv0d0 U5802 ( .I(dbg_uart_wishbone_dat_w[27]), .ZN(n5471) );
  inv0d0 U5803 ( .I(mgmtsoc_ibus_ibus_dat_r[27]), .ZN(n5470) );
  oai222d1 U5804 ( .A1(n5481), .A2(n5471), .B1(n5485), .B2(n5470), .C1(n5469), 
        .C2(n5482), .ZN(n3256) );
  inv0d0 U5805 ( .I(dbg_uart_wishbone_dat_w[28]), .ZN(n5474) );
  inv0d0 U5806 ( .I(mgmtsoc_ibus_ibus_dat_r[28]), .ZN(n5473) );
  oai222d1 U5807 ( .A1(n5487), .A2(n5474), .B1(n5485), .B2(n5473), .C1(n5472), 
        .C2(n5482), .ZN(n3255) );
  inv0d0 U5808 ( .I(dbg_uart_wishbone_dat_w[29]), .ZN(n5477) );
  inv0d0 U5809 ( .I(mgmtsoc_ibus_ibus_dat_r[29]), .ZN(n5476) );
  oai222d1 U5810 ( .A1(n5487), .A2(n5477), .B1(n5485), .B2(n5476), .C1(n5475), 
        .C2(n5482), .ZN(n3254) );
  inv0d0 U5811 ( .I(dbg_uart_wishbone_dat_w[30]), .ZN(n5480) );
  inv0d0 U5812 ( .I(mgmtsoc_ibus_ibus_dat_r[30]), .ZN(n5479) );
  oai222d1 U5813 ( .A1(n5481), .A2(n5480), .B1(n5485), .B2(n5479), .C1(n5478), 
        .C2(n5482), .ZN(n3253) );
  inv0d0 U5814 ( .I(dbg_uart_wishbone_dat_w[31]), .ZN(n5486) );
  inv0d0 U5815 ( .I(mgmtsoc_ibus_ibus_dat_r[31]), .ZN(n5484) );
  oai222d1 U5816 ( .A1(n5487), .A2(n5486), .B1(n5485), .B2(n5484), .C1(n5483), 
        .C2(n5482), .ZN(n3252) );
  nd04d1 U5817 ( .A1(n5490), .A2(n5489), .A3(N5758), .A4(n5488), .ZN(n5599) );
  inv0d1 U5818 ( .I(n5599), .ZN(n5605) );
  nr03d1 U5819 ( .A1(n5492), .A2(n5605), .A3(n5491), .ZN(n5519) );
  aoi22d1 U5820 ( .A1(dbg_uart_wishbone_adr[0]), .A2(n5519), .B1(n5604), .B2(
        n5493), .ZN(n5494) );
  oai21d1 U5821 ( .B1(n5969), .B2(n5599), .A(n5494), .ZN(n3251) );
  buffd1 U5822 ( .I(n5592), .Z(n5571) );
  ah01d1 U5823 ( .A(dbg_uart_wishbone_adr[0]), .B(dbg_uart_incr), .CO(n5497), 
        .S(n5493) );
  aoi22d1 U5824 ( .A1(dbg_uart_wishbone_adr[1]), .A2(n5519), .B1(n5571), .B2(
        n5495), .ZN(n5496) );
  oai21d1 U5825 ( .B1(n5970), .B2(n5599), .A(n5496), .ZN(n3250) );
  ah01d1 U5826 ( .A(n5497), .B(dbg_uart_wishbone_adr[1]), .CO(n5500), .S(n5495) );
  aoi22d1 U5827 ( .A1(dbg_uart_wishbone_adr[2]), .A2(n5519), .B1(n5571), .B2(
        n5498), .ZN(n5499) );
  oai21d1 U5828 ( .B1(n5971), .B2(n5599), .A(n5499), .ZN(n3249) );
  ah01d1 U5829 ( .A(n5500), .B(dbg_uart_wishbone_adr[2]), .CO(n5503), .S(n5498) );
  aoi22d1 U5830 ( .A1(dbg_uart_wishbone_adr[3]), .A2(n5519), .B1(n5571), .B2(
        n5501), .ZN(n5502) );
  oai21d1 U5831 ( .B1(n5972), .B2(n5599), .A(n5502), .ZN(n3248) );
  ah01d1 U5832 ( .A(n5503), .B(dbg_uart_wishbone_adr[3]), .CO(n5506), .S(n5501) );
  aoi22d1 U5833 ( .A1(dbg_uart_wishbone_adr[4]), .A2(n5519), .B1(n5571), .B2(
        n5504), .ZN(n5505) );
  oai21d1 U5834 ( .B1(n5973), .B2(n5599), .A(n5505), .ZN(n3247) );
  ah01d1 U5835 ( .A(n5506), .B(dbg_uart_wishbone_adr[4]), .CO(n5509), .S(n5504) );
  aoi22d1 U5836 ( .A1(dbg_uart_wishbone_adr[5]), .A2(n5519), .B1(n5571), .B2(
        n5507), .ZN(n5508) );
  oai21d1 U5837 ( .B1(n5974), .B2(n5599), .A(n5508), .ZN(n3246) );
  ah01d1 U5838 ( .A(n5509), .B(dbg_uart_wishbone_adr[5]), .CO(n5512), .S(n5507) );
  aoi22d1 U5839 ( .A1(dbg_uart_wishbone_adr[6]), .A2(n5519), .B1(n5571), .B2(
        n5510), .ZN(n5511) );
  oai21d1 U5840 ( .B1(n5975), .B2(n5599), .A(n5511), .ZN(n3245) );
  ah01d1 U5841 ( .A(n5512), .B(dbg_uart_wishbone_adr[6]), .CO(n5515), .S(n5510) );
  aoi22d1 U5842 ( .A1(dbg_uart_wishbone_adr[7]), .A2(n5519), .B1(n5571), .B2(
        n5513), .ZN(n5514) );
  oai21d1 U5843 ( .B1(n5976), .B2(n5599), .A(n5514), .ZN(n3244) );
  ah01d1 U5844 ( .A(n5515), .B(dbg_uart_wishbone_adr[7]), .CO(n5520), .S(n5513) );
  aoi22d1 U5845 ( .A1(dbg_uart_wishbone_adr[8]), .A2(n5519), .B1(n5571), .B2(
        n5516), .ZN(n5517) );
  oai21d1 U5846 ( .B1(n5518), .B2(n5599), .A(n5517), .ZN(n3243) );
  buffd1 U5847 ( .I(n5519), .Z(n5597) );
  ah01d1 U5848 ( .A(n5520), .B(dbg_uart_wishbone_adr[8]), .CO(n5524), .S(n5516) );
  aoi22d1 U5849 ( .A1(dbg_uart_wishbone_adr[9]), .A2(n5597), .B1(n5571), .B2(
        n5521), .ZN(n5522) );
  oai21d1 U5850 ( .B1(n5523), .B2(n5599), .A(n5522), .ZN(n3242) );
  ah01d1 U5851 ( .A(n5524), .B(dbg_uart_wishbone_adr[9]), .CO(n5528), .S(n5521) );
  aoi22d1 U5852 ( .A1(dbg_uart_wishbone_adr[10]), .A2(n5597), .B1(n5571), .B2(
        n5525), .ZN(n5526) );
  oai21d1 U5853 ( .B1(n5527), .B2(n5599), .A(n5526), .ZN(n3241) );
  inv0d1 U5854 ( .I(n5597), .ZN(n5607) );
  ah01d1 U5855 ( .A(n5528), .B(dbg_uart_wishbone_adr[10]), .CO(n5531), .S(
        n5525) );
  aoi22d1 U5856 ( .A1(dbg_uart_wishbone_adr[3]), .A2(n5605), .B1(n5571), .B2(
        n5529), .ZN(n5530) );
  oai21d1 U5857 ( .B1(n5561), .B2(n5607), .A(n5530), .ZN(n3240) );
  ah01d1 U5858 ( .A(n5531), .B(dbg_uart_wishbone_adr[11]), .CO(n5535), .S(
        n5529) );
  aoi22d1 U5859 ( .A1(dbg_uart_wishbone_adr[4]), .A2(n5605), .B1(n5571), .B2(
        n5532), .ZN(n5533) );
  oai21d1 U5860 ( .B1(n5534), .B2(n5607), .A(n5533), .ZN(n3239) );
  ah01d1 U5861 ( .A(n5535), .B(dbg_uart_wishbone_adr[12]), .CO(n5538), .S(
        n5532) );
  aoi22d1 U5862 ( .A1(dbg_uart_wishbone_adr[5]), .A2(n5605), .B1(n5604), .B2(
        n5536), .ZN(n5537) );
  oai21d1 U5863 ( .B1(n5568), .B2(n5607), .A(n5537), .ZN(n3238) );
  ah01d1 U5864 ( .A(n5538), .B(dbg_uart_wishbone_adr[13]), .CO(n5542), .S(
        n5536) );
  aoi22d1 U5865 ( .A1(dbg_uart_wishbone_adr[14]), .A2(n5597), .B1(n5604), .B2(
        n5539), .ZN(n5540) );
  oai21d1 U5866 ( .B1(n5541), .B2(n5599), .A(n5540), .ZN(n3237) );
  ah01d1 U5867 ( .A(n5542), .B(dbg_uart_wishbone_adr[14]), .CO(n5546), .S(
        n5539) );
  aoi22d1 U5868 ( .A1(dbg_uart_wishbone_adr[7]), .A2(n5605), .B1(n5604), .B2(
        n5543), .ZN(n5544) );
  oai21d1 U5869 ( .B1(n5545), .B2(n5607), .A(n5544), .ZN(n3236) );
  ah01d1 U5870 ( .A(n5546), .B(dbg_uart_wishbone_adr[15]), .CO(n5550), .S(
        n5543) );
  aoi22d1 U5871 ( .A1(dbg_uart_wishbone_adr[8]), .A2(n5605), .B1(n5571), .B2(
        n5547), .ZN(n5548) );
  oai21d1 U5872 ( .B1(n5549), .B2(n5607), .A(n5548), .ZN(n3235) );
  ah01d1 U5873 ( .A(n5550), .B(dbg_uart_wishbone_adr[16]), .CO(n5554), .S(
        n5547) );
  aoi22d1 U5874 ( .A1(dbg_uart_wishbone_adr[9]), .A2(n5605), .B1(n5604), .B2(
        n5551), .ZN(n5552) );
  oai21d1 U5875 ( .B1(n5553), .B2(n5607), .A(n5552), .ZN(n3234) );
  ah01d1 U5876 ( .A(n5554), .B(dbg_uart_wishbone_adr[17]), .CO(n5558), .S(
        n5551) );
  aoi22d1 U5877 ( .A1(dbg_uart_wishbone_adr[10]), .A2(n5605), .B1(n5571), .B2(
        n5555), .ZN(n5556) );
  oai21d1 U5878 ( .B1(n5557), .B2(n5607), .A(n5556), .ZN(n3233) );
  ah01d1 U5879 ( .A(n5558), .B(dbg_uart_wishbone_adr[18]), .CO(n5562), .S(
        n5555) );
  aoi22d1 U5880 ( .A1(dbg_uart_wishbone_adr[19]), .A2(n5597), .B1(n5592), .B2(
        n5559), .ZN(n5560) );
  oai21d1 U5881 ( .B1(n5561), .B2(n5599), .A(n5560), .ZN(n3232) );
  ah01d1 U5882 ( .A(n5562), .B(dbg_uart_wishbone_adr[19]), .CO(n5565), .S(
        n5559) );
  aoi22d1 U5883 ( .A1(dbg_uart_wishbone_adr[12]), .A2(n5605), .B1(n5604), .B2(
        n5563), .ZN(n5564) );
  oai21d1 U5884 ( .B1(n5600), .B2(n5607), .A(n5564), .ZN(n3231) );
  ah01d1 U5885 ( .A(n5565), .B(dbg_uart_wishbone_adr[20]), .CO(n5569), .S(
        n5563) );
  aoi22d1 U5886 ( .A1(dbg_uart_wishbone_adr[21]), .A2(n5597), .B1(n5571), .B2(
        n5566), .ZN(n5567) );
  oai21d1 U5887 ( .B1(n5568), .B2(n5599), .A(n5567), .ZN(n3230) );
  ah01d1 U5888 ( .A(n5569), .B(dbg_uart_wishbone_adr[21]), .CO(n5574), .S(
        n5566) );
  aoi22d1 U5889 ( .A1(dbg_uart_wishbone_adr[14]), .A2(n5605), .B1(n5571), .B2(
        n5570), .ZN(n5572) );
  oai21d1 U5890 ( .B1(n5573), .B2(n5607), .A(n5572), .ZN(n3229) );
  ah01d1 U5891 ( .A(n5574), .B(dbg_uart_wishbone_adr[22]), .CO(n5578), .S(
        n5570) );
  aoi22d1 U5892 ( .A1(dbg_uart_wishbone_adr[15]), .A2(n5605), .B1(n5604), .B2(
        n5575), .ZN(n5576) );
  oai21d1 U5893 ( .B1(n5577), .B2(n5607), .A(n5576), .ZN(n3228) );
  ah01d1 U5894 ( .A(n5578), .B(dbg_uart_wishbone_adr[23]), .CO(n5582), .S(
        n5575) );
  aoi22d1 U5895 ( .A1(dbg_uart_wishbone_adr[16]), .A2(n5605), .B1(n5592), .B2(
        n5579), .ZN(n5580) );
  oai21d1 U5896 ( .B1(n5581), .B2(n5607), .A(n5580), .ZN(n3227) );
  ah01d1 U5897 ( .A(n5582), .B(dbg_uart_wishbone_adr[24]), .CO(n5586), .S(
        n5579) );
  aoi22d1 U5898 ( .A1(dbg_uart_wishbone_adr[17]), .A2(n5605), .B1(n5592), .B2(
        n5583), .ZN(n5584) );
  oai21d1 U5899 ( .B1(n5585), .B2(n5607), .A(n5584), .ZN(n3226) );
  ah01d1 U5900 ( .A(n5586), .B(dbg_uart_wishbone_adr[25]), .CO(n5590), .S(
        n5583) );
  aoi22d1 U5901 ( .A1(dbg_uart_wishbone_adr[18]), .A2(n5605), .B1(n5592), .B2(
        n5587), .ZN(n5588) );
  oai21d1 U5902 ( .B1(n5589), .B2(n5607), .A(n5588), .ZN(n3225) );
  ah01d1 U5903 ( .A(n5590), .B(dbg_uart_wishbone_adr[26]), .CO(n5595), .S(
        n5587) );
  aoi22d1 U5904 ( .A1(dbg_uart_wishbone_adr[19]), .A2(n5605), .B1(n5592), .B2(
        n5591), .ZN(n5593) );
  oai21d1 U5905 ( .B1(n5594), .B2(n5607), .A(n5593), .ZN(n3224) );
  ah01d1 U5906 ( .A(n5595), .B(dbg_uart_wishbone_adr[27]), .CO(n5601), .S(
        n5591) );
  aoi22d1 U5907 ( .A1(dbg_uart_wishbone_adr[28]), .A2(n5597), .B1(n5604), .B2(
        n5596), .ZN(n5598) );
  oai21d1 U5908 ( .B1(n5600), .B2(n5599), .A(n5598), .ZN(n3223) );
  ah01d1 U5909 ( .A(n5601), .B(dbg_uart_wishbone_adr[28]), .CO(n5602), .S(
        n5596) );
  ah01d1 U5910 ( .A(n5602), .B(dbg_uart_wishbone_adr[29]), .S(n5603) );
  aoi22d1 U5911 ( .A1(dbg_uart_wishbone_adr[21]), .A2(n5605), .B1(n5604), .B2(
        n5603), .ZN(n5606) );
  oai21d1 U5912 ( .B1(n5608), .B2(n5607), .A(n5606), .ZN(n3222) );
  nr02d1 U5913 ( .A1(n5664), .A2(n5707), .ZN(n5727) );
  buffd1 U5914 ( .I(n5727), .Z(n5710) );
  aoi22d1 U5915 ( .A1(mgmtsoc_litespimmap_burst_adr[0]), .A2(n5710), .B1(n5664), .B2(n5609), .ZN(n5610) );
  oai21d1 U5916 ( .B1(n5611), .B2(n5721), .A(n5610), .ZN(n3221) );
  aoi22d1 U5917 ( .A1(mgmtsoc_litespimmap_burst_adr[1]), .A2(n5710), .B1(n5664), .B2(n5612), .ZN(n5613) );
  oai21d1 U5918 ( .B1(n5614), .B2(n5721), .A(n5613), .ZN(n3220) );
  ah01d1 U5919 ( .A(mgmtsoc_litespimmap_burst_adr[0]), .B(
        mgmtsoc_litespimmap_burst_adr[1]), .CO(n5618), .S(n5612) );
  aoi22d1 U5920 ( .A1(mgmtsoc_litespimmap_burst_adr[2]), .A2(n5710), .B1(n5664), .B2(n5615), .ZN(n5616) );
  oai21d1 U5921 ( .B1(n5617), .B2(n5721), .A(n5616), .ZN(n3219) );
  ah01d1 U5922 ( .A(n5618), .B(mgmtsoc_litespimmap_burst_adr[2]), .CO(n5622), 
        .S(n5615) );
  aoi22d1 U5923 ( .A1(mgmtsoc_litespimmap_burst_adr[3]), .A2(n5710), .B1(n5664), .B2(n5619), .ZN(n5620) );
  oai21d1 U5924 ( .B1(n5621), .B2(n5721), .A(n5620), .ZN(n3218) );
  ah01d1 U5925 ( .A(n5622), .B(mgmtsoc_litespimmap_burst_adr[3]), .CO(n5626), 
        .S(n5619) );
  aoi22d1 U5926 ( .A1(mgmtsoc_litespimmap_burst_adr[4]), .A2(n5710), .B1(n5664), .B2(n5623), .ZN(n5624) );
  oai21d1 U5927 ( .B1(n5625), .B2(n5721), .A(n5624), .ZN(n3217) );
  buffd1 U5928 ( .I(n5726), .Z(n5719) );
  ah01d1 U5929 ( .A(n5626), .B(mgmtsoc_litespimmap_burst_adr[4]), .CO(n5630), 
        .S(n5623) );
  aoi22d1 U5930 ( .A1(mgmtsoc_litespimmap_burst_adr[5]), .A2(n5710), .B1(n5719), .B2(n5627), .ZN(n5628) );
  oai21d1 U5931 ( .B1(n5629), .B2(n5721), .A(n5628), .ZN(n3216) );
  ah01d1 U5932 ( .A(n5630), .B(mgmtsoc_litespimmap_burst_adr[5]), .CO(n5634), 
        .S(n5627) );
  aoi22d1 U5933 ( .A1(mgmtsoc_litespimmap_burst_adr[6]), .A2(n5710), .B1(n5726), .B2(n5631), .ZN(n5632) );
  oai21d1 U5934 ( .B1(n5633), .B2(n5721), .A(n5632), .ZN(n3215) );
  ah01d1 U5935 ( .A(n5634), .B(mgmtsoc_litespimmap_burst_adr[6]), .CO(n5638), 
        .S(n5631) );
  aoi22d1 U5936 ( .A1(mgmtsoc_litespimmap_burst_adr[7]), .A2(n5710), .B1(n5726), .B2(n5635), .ZN(n5636) );
  oai21d1 U5937 ( .B1(n5637), .B2(n5721), .A(n5636), .ZN(n3214) );
  ah01d1 U5938 ( .A(n5638), .B(mgmtsoc_litespimmap_burst_adr[7]), .CO(n5642), 
        .S(n5635) );
  aoi22d1 U5939 ( .A1(mgmtsoc_litespimmap_burst_adr[8]), .A2(n5710), .B1(n5664), .B2(n5639), .ZN(n5640) );
  oai21d1 U5940 ( .B1(n5641), .B2(n5729), .A(n5640), .ZN(n3213) );
  ah01d1 U5941 ( .A(n5642), .B(mgmtsoc_litespimmap_burst_adr[8]), .CO(n5646), 
        .S(n5639) );
  aoi22d1 U5942 ( .A1(mgmtsoc_litespimmap_burst_adr[9]), .A2(n5727), .B1(n5664), .B2(n5643), .ZN(n5644) );
  oai21d1 U5943 ( .B1(n5645), .B2(n5721), .A(n5644), .ZN(n3212) );
  ah01d1 U5944 ( .A(n5646), .B(mgmtsoc_litespimmap_burst_adr[9]), .CO(n5650), 
        .S(n5643) );
  aoi22d1 U5945 ( .A1(mgmtsoc_litespimmap_burst_adr[10]), .A2(n5710), .B1(
        n5719), .B2(n5647), .ZN(n5648) );
  oai21d1 U5946 ( .B1(n5649), .B2(n5721), .A(n5648), .ZN(n3211) );
  ah01d1 U5947 ( .A(n5650), .B(mgmtsoc_litespimmap_burst_adr[10]), .CO(n5654), 
        .S(n5647) );
  aoi22d1 U5948 ( .A1(mgmtsoc_litespimmap_burst_adr[11]), .A2(n5710), .B1(
        n5719), .B2(n5651), .ZN(n5652) );
  oai21d1 U5949 ( .B1(n5653), .B2(n5721), .A(n5652), .ZN(n3210) );
  ah01d1 U5950 ( .A(n5654), .B(mgmtsoc_litespimmap_burst_adr[11]), .CO(n5658), 
        .S(n5651) );
  aoi22d1 U5951 ( .A1(mgmtsoc_litespimmap_burst_adr[12]), .A2(n5727), .B1(
        n5719), .B2(n5655), .ZN(n5656) );
  oai21d1 U5952 ( .B1(n5657), .B2(n5721), .A(n5656), .ZN(n3209) );
  ah01d1 U5953 ( .A(n5658), .B(mgmtsoc_litespimmap_burst_adr[12]), .CO(n5662), 
        .S(n5655) );
  aoi22d1 U5954 ( .A1(mgmtsoc_litespimmap_burst_adr[13]), .A2(n5727), .B1(
        n5719), .B2(n5659), .ZN(n5660) );
  oai21d1 U5955 ( .B1(n5661), .B2(n5721), .A(n5660), .ZN(n3208) );
  ah01d1 U5956 ( .A(n5662), .B(mgmtsoc_litespimmap_burst_adr[13]), .CO(n5667), 
        .S(n5659) );
  aoi22d1 U5957 ( .A1(mgmtsoc_litespimmap_burst_adr[14]), .A2(n5727), .B1(
        n5664), .B2(n5663), .ZN(n5665) );
  oai21d1 U5958 ( .B1(n5666), .B2(n5721), .A(n5665), .ZN(n3207) );
  ah01d1 U5959 ( .A(n5667), .B(mgmtsoc_litespimmap_burst_adr[14]), .CO(n5671), 
        .S(n5663) );
  aoi22d1 U5960 ( .A1(mgmtsoc_litespimmap_burst_adr[15]), .A2(n5710), .B1(
        n5719), .B2(n5668), .ZN(n5669) );
  oai21d1 U5961 ( .B1(n5670), .B2(n5721), .A(n5669), .ZN(n3206) );
  ah01d1 U5962 ( .A(n5671), .B(mgmtsoc_litespimmap_burst_adr[15]), .CO(n5675), 
        .S(n5668) );
  aoi22d1 U5963 ( .A1(mgmtsoc_litespimmap_burst_adr[16]), .A2(n5710), .B1(
        n5719), .B2(n5672), .ZN(n5673) );
  oai21d1 U5964 ( .B1(n5674), .B2(n5721), .A(n5673), .ZN(n3205) );
  ah01d1 U5965 ( .A(n5675), .B(mgmtsoc_litespimmap_burst_adr[16]), .CO(n5679), 
        .S(n5672) );
  aoi22d1 U5966 ( .A1(mgmtsoc_litespimmap_burst_adr[17]), .A2(n5710), .B1(
        n5726), .B2(n5676), .ZN(n5677) );
  oai21d1 U5967 ( .B1(n5678), .B2(n5721), .A(n5677), .ZN(n3204) );
  ah01d1 U5968 ( .A(n5679), .B(mgmtsoc_litespimmap_burst_adr[17]), .CO(n5683), 
        .S(n5676) );
  aoi22d1 U5969 ( .A1(mgmtsoc_litespimmap_burst_adr[18]), .A2(n5710), .B1(
        n5719), .B2(n5680), .ZN(n5681) );
  oai21d1 U5970 ( .B1(n5682), .B2(n5721), .A(n5681), .ZN(n3203) );
  ah01d1 U5971 ( .A(n5683), .B(mgmtsoc_litespimmap_burst_adr[18]), .CO(n5687), 
        .S(n5680) );
  aoi22d1 U5972 ( .A1(mgmtsoc_litespimmap_burst_adr[19]), .A2(n5727), .B1(
        n5726), .B2(n5684), .ZN(n5685) );
  oai21d1 U5973 ( .B1(n5686), .B2(n5721), .A(n5685), .ZN(n3202) );
  ah01d1 U5974 ( .A(n5687), .B(mgmtsoc_litespimmap_burst_adr[19]), .CO(n5691), 
        .S(n5684) );
  aoi22d1 U5975 ( .A1(mgmtsoc_litespimmap_burst_adr[20]), .A2(n5710), .B1(
        n5719), .B2(n5688), .ZN(n5689) );
  oai21d1 U5976 ( .B1(n5690), .B2(n5721), .A(n5689), .ZN(n3201) );
  ah01d1 U5977 ( .A(n5691), .B(mgmtsoc_litespimmap_burst_adr[20]), .CO(n5695), 
        .S(n5688) );
  aoi22d1 U5978 ( .A1(mgmtsoc_litespimmap_burst_adr[21]), .A2(n5727), .B1(
        n5719), .B2(n5692), .ZN(n5693) );
  oai21d1 U5979 ( .B1(n5694), .B2(n5721), .A(n5693), .ZN(n3200) );
  ah01d1 U5980 ( .A(n5695), .B(mgmtsoc_litespimmap_burst_adr[21]), .CO(n5698), 
        .S(n5692) );
  aoi22d1 U5981 ( .A1(mgmtsoc_litespimmap_burst_adr[22]), .A2(n5727), .B1(
        n5719), .B2(n5696), .ZN(n5697) );
  oaim21d1 U5982 ( .B1(mprj_adr_o[24]), .B2(n5707), .A(n5697), .ZN(n3199) );
  ah01d1 U5983 ( .A(n5698), .B(mgmtsoc_litespimmap_burst_adr[22]), .CO(n5701), 
        .S(n5696) );
  aoi22d1 U5984 ( .A1(mgmtsoc_litespimmap_burst_adr[23]), .A2(n5727), .B1(
        n5719), .B2(n5699), .ZN(n5700) );
  oaim21d1 U5985 ( .B1(mprj_adr_o[25]), .B2(n5707), .A(n5700), .ZN(n3198) );
  ah01d1 U5986 ( .A(n5701), .B(mgmtsoc_litespimmap_burst_adr[23]), .CO(n5704), 
        .S(n5699) );
  aoi22d1 U5987 ( .A1(mgmtsoc_litespimmap_burst_adr[24]), .A2(n5727), .B1(
        n5719), .B2(n5702), .ZN(n5703) );
  oaim21d1 U5988 ( .B1(mprj_adr_o[26]), .B2(n5707), .A(n5703), .ZN(n3197) );
  ah01d1 U5989 ( .A(n5704), .B(mgmtsoc_litespimmap_burst_adr[24]), .CO(n5708), 
        .S(n5702) );
  aoi22d1 U5990 ( .A1(mgmtsoc_litespimmap_burst_adr[25]), .A2(n5727), .B1(
        n5719), .B2(n5705), .ZN(n5706) );
  oaim21d1 U5991 ( .B1(mprj_adr_o[27]), .B2(n5707), .A(n5706), .ZN(n3196) );
  ah01d1 U5992 ( .A(n5708), .B(mgmtsoc_litespimmap_burst_adr[25]), .CO(n5713), 
        .S(n5705) );
  aoi22d1 U5993 ( .A1(mgmtsoc_litespimmap_burst_adr[26]), .A2(n5710), .B1(
        n5719), .B2(n5709), .ZN(n5711) );
  oai21d1 U5994 ( .B1(n5712), .B2(n5721), .A(n5711), .ZN(n3195) );
  ah01d1 U5995 ( .A(n5713), .B(mgmtsoc_litespimmap_burst_adr[26]), .CO(n5717), 
        .S(n5709) );
  aoi22d1 U5996 ( .A1(mgmtsoc_litespimmap_burst_adr[27]), .A2(n5727), .B1(
        n5719), .B2(n5714), .ZN(n5715) );
  oai21d1 U5997 ( .B1(n5716), .B2(n5721), .A(n5715), .ZN(n3194) );
  ah01d1 U5998 ( .A(n5717), .B(mgmtsoc_litespimmap_burst_adr[27]), .CO(n5723), 
        .S(n5714) );
  aoi22d1 U5999 ( .A1(mgmtsoc_litespimmap_burst_adr[28]), .A2(n5727), .B1(
        n5719), .B2(n5718), .ZN(n5720) );
  oai21d1 U6000 ( .B1(n5722), .B2(n5721), .A(n5720), .ZN(n3193) );
  ah01d1 U6001 ( .A(n5723), .B(mgmtsoc_litespimmap_burst_adr[28]), .CO(n5724), 
        .S(n5718) );
  xr02d1 U6002 ( .A1(n5724), .A2(mgmtsoc_litespimmap_burst_adr[29]), .Z(n5725)
         );
  aoi22d1 U6003 ( .A1(mgmtsoc_litespimmap_burst_adr[29]), .A2(n5727), .B1(
        n5726), .B2(n5725), .ZN(n5728) );
  oai21d1 U6004 ( .B1(n5730), .B2(n5729), .A(n5728), .ZN(n3192) );
  inv0d0 U6005 ( .I(mgmtsoc_litespisdrphycore_posedge_reg2), .ZN(n5731) );
  oan211d1 U6006 ( .C1(n5734), .C2(n5733), .B(n5732), .A(n5731), .ZN(n5737) );
  nd02d1 U6007 ( .A1(n5737), .A2(n5735), .ZN(n5774) );
  buffd1 U6008 ( .I(n5774), .Z(n5765) );
  nd02d1 U6009 ( .A1(n5737), .A2(n5736), .ZN(n5768) );
  buffd1 U6010 ( .I(n5768), .Z(n5772) );
  nd02d1 U6011 ( .A1(n5765), .A2(n5772), .ZN(n5776) );
  oai222d1 U6012 ( .A1(n5776), .A2(n5771), .B1(n5765), .B2(n5767), .C1(n5772), 
        .C2(n5773), .ZN(n3191) );
  buffd1 U6013 ( .I(n5776), .Z(n5770) );
  inv0d0 U6014 ( .I(\mgmtsoc_litespisdrphycore_dq_i[1] ), .ZN(n5738) );
  oai22d1 U6015 ( .A1(n5739), .A2(n5770), .B1(n5772), .B2(n5738), .ZN(n3190)
         );
  oai222d1 U6016 ( .A1(n5738), .A2(n5765), .B1(n5772), .B2(n5739), .C1(n5770), 
        .C2(n5740), .ZN(n3189) );
  oai222d1 U6017 ( .A1(n5770), .A2(n5741), .B1(n5765), .B2(n5739), .C1(n5772), 
        .C2(n5740), .ZN(n3188) );
  oai222d1 U6018 ( .A1(n5770), .A2(n5742), .B1(n5765), .B2(n5740), .C1(n5772), 
        .C2(n5741), .ZN(n3187) );
  oai222d1 U6019 ( .A1(n5770), .A2(n5743), .B1(n5765), .B2(n5741), .C1(n5768), 
        .C2(n5742), .ZN(n3186) );
  oai222d1 U6020 ( .A1(n5770), .A2(n5744), .B1(n5774), .B2(n5742), .C1(n5768), 
        .C2(n5743), .ZN(n3185) );
  oai222d1 U6021 ( .A1(n5770), .A2(n5745), .B1(n5765), .B2(n5743), .C1(n5768), 
        .C2(n5744), .ZN(n3184) );
  oai222d1 U6022 ( .A1(n5776), .A2(n5746), .B1(n5765), .B2(n5744), .C1(n5768), 
        .C2(n5745), .ZN(n3183) );
  oai222d1 U6023 ( .A1(n5770), .A2(n5747), .B1(n5774), .B2(n5745), .C1(n5768), 
        .C2(n5746), .ZN(n3182) );
  oai222d1 U6024 ( .A1(n5776), .A2(n5748), .B1(n5765), .B2(n5746), .C1(n5768), 
        .C2(n5747), .ZN(n3181) );
  oai222d1 U6025 ( .A1(n5770), .A2(n5749), .B1(n5774), .B2(n5747), .C1(n5768), 
        .C2(n5748), .ZN(n3180) );
  oai222d1 U6026 ( .A1(n5770), .A2(n5750), .B1(n5774), .B2(n5748), .C1(n5768), 
        .C2(n5749), .ZN(n3179) );
  oai222d1 U6027 ( .A1(n5770), .A2(n5751), .B1(n5774), .B2(n5749), .C1(n5768), 
        .C2(n5750), .ZN(n3178) );
  oai222d1 U6028 ( .A1(n5776), .A2(n5752), .B1(n5765), .B2(n5750), .C1(n5772), 
        .C2(n5751), .ZN(n3177) );
  oai222d1 U6029 ( .A1(n5770), .A2(n5753), .B1(n5765), .B2(n5751), .C1(n5768), 
        .C2(n5752), .ZN(n3176) );
  oai222d1 U6030 ( .A1(n5770), .A2(n5754), .B1(n5765), .B2(n5752), .C1(n5768), 
        .C2(n5753), .ZN(n3175) );
  oai222d1 U6031 ( .A1(n5776), .A2(n5755), .B1(n5765), .B2(n5753), .C1(n5768), 
        .C2(n5754), .ZN(n3174) );
  oai222d1 U6032 ( .A1(n5770), .A2(n5756), .B1(n5774), .B2(n5754), .C1(n5772), 
        .C2(n5755), .ZN(n3173) );
  oai222d1 U6033 ( .A1(n5776), .A2(n5757), .B1(n5774), .B2(n5755), .C1(n5772), 
        .C2(n5756), .ZN(n3172) );
  oai222d1 U6034 ( .A1(n5776), .A2(n5758), .B1(n5774), .B2(n5756), .C1(n5772), 
        .C2(n5757), .ZN(n3171) );
  oai222d1 U6035 ( .A1(n5770), .A2(n5759), .B1(n5774), .B2(n5757), .C1(n5772), 
        .C2(n5758), .ZN(n3170) );
  oai222d1 U6036 ( .A1(n5776), .A2(n5760), .B1(n5765), .B2(n5758), .C1(n5772), 
        .C2(n5759), .ZN(n3169) );
  oai222d1 U6037 ( .A1(n5776), .A2(n5761), .B1(n5774), .B2(n5759), .C1(n5772), 
        .C2(n5760), .ZN(n3168) );
  oai222d1 U6038 ( .A1(n5776), .A2(n5762), .B1(n5765), .B2(n5760), .C1(n5768), 
        .C2(n5761), .ZN(n3167) );
  oai222d1 U6039 ( .A1(n5776), .A2(n5763), .B1(n5774), .B2(n5761), .C1(n5768), 
        .C2(n5762), .ZN(n3166) );
  oai222d1 U6040 ( .A1(n5776), .A2(n5764), .B1(n5774), .B2(n5762), .C1(n5772), 
        .C2(n5763), .ZN(n3165) );
  oai222d1 U6041 ( .A1(n5776), .A2(n5766), .B1(n5765), .B2(n5763), .C1(n5772), 
        .C2(n5764), .ZN(n3164) );
  oai222d1 U6042 ( .A1(n5770), .A2(n5769), .B1(n5765), .B2(n5764), .C1(n5768), 
        .C2(n5766), .ZN(n3163) );
  oai222d1 U6043 ( .A1(n5776), .A2(n5767), .B1(n5774), .B2(n5766), .C1(n5772), 
        .C2(n5769), .ZN(n3162) );
  oai222d1 U6044 ( .A1(n5770), .A2(n5773), .B1(n5774), .B2(n5769), .C1(n5768), 
        .C2(n5767), .ZN(n3161) );
  oai222d1 U6045 ( .A1(n5776), .A2(n5775), .B1(n5774), .B2(n5773), .C1(n5772), 
        .C2(n5771), .ZN(n3160) );
  inv0d0 U6046 ( .I(mgmtsoc_litespisdrphycore_sr_out[0]), .ZN(n5909) );
  inv0d0 U6047 ( .I(n5777), .ZN(n5779) );
  nr02d0 U6048 ( .A1(n5779), .A2(n5778), .ZN(n5880) );
  oaim22d1 U6049 ( .A1(n5906), .A2(n5909), .B1(n5780), .B2(n5880), .ZN(n3159)
         );
  an02d0 U6050 ( .A1(n5784), .A2(n5785), .Z(n5881) );
  aoi22d1 U6051 ( .A1(n5893), .A2(mgmtsoc_litespisdrphycore_sr_out[27]), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[23]), .ZN(n5782) );
  aoi22d1 U6052 ( .A1(n5871), .A2(mgmtsoc_litespisdrphycore_sr_out[31]), .B1(
        n5886), .B2(mgmtsoc_litespisdrphycore_sr_out[29]), .ZN(n5781) );
  oai211d1 U6053 ( .C1(n5908), .C2(n5799), .A(n5782), .B(n5781), .ZN(n5795) );
  or02d1 U6054 ( .A1(n5786), .A2(n5785), .Z(n5910) );
  aoi22d1 U6055 ( .A1(n5787), .A2(
        mgmtsoc_port_master_user_port_sink_payload_data[28]), .B1(n5789), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[29]), .ZN(n5816) );
  aoi22d1 U6056 ( .A1(n5787), .A2(
        mgmtsoc_port_master_user_port_sink_payload_data[30]), .B1(n5800), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[31]), .ZN(n5788) );
  aoi22d1 U6057 ( .A1(n5790), .A2(n5816), .B1(n5788), .B2(n5804), .ZN(n5791)
         );
  aoi22d1 U6058 ( .A1(n5801), .A2(
        mgmtsoc_port_master_user_port_sink_payload_data[24]), .B1(n5789), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[25]), .ZN(n5819) );
  aoi22d1 U6059 ( .A1(n5801), .A2(
        mgmtsoc_port_master_user_port_sink_payload_data[26]), .B1(n5800), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[27]), .ZN(n5817) );
  aoi22d1 U6060 ( .A1(n5790), .A2(n5819), .B1(n5817), .B2(n5804), .ZN(n5832)
         );
  aoi22d1 U6061 ( .A1(n5862), .A2(n5791), .B1(n5832), .B2(n5830), .ZN(n5792)
         );
  oai22d1 U6062 ( .A1(n5877), .A2(n5793), .B1(n5910), .B2(n5792), .ZN(n5794)
         );
  aor211d1 U6063 ( .C1(n5881), .C2(n5796), .A(n5795), .B(n5794), .Z(n3158) );
  aoi22d1 U6064 ( .A1(mgmtsoc_litespisdrphycore_sr_out[26]), .A2(n5885), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[22]), .ZN(n5798) );
  aoi22d1 U6065 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[29]), .B1(
        mgmtsoc_litespisdrphycore_sr_out[28]), .B2(n5886), .ZN(n5797) );
  oai211d1 U6066 ( .C1(n5906), .C2(n5799), .A(n5798), .B(n5797), .ZN(n5811) );
  aoi22d1 U6067 ( .A1(n5801), .A2(
        mgmtsoc_port_master_user_port_sink_payload_data[29]), .B1(n5800), .B2(
        mgmtsoc_port_master_user_port_sink_payload_data[30]), .ZN(n5802) );
  aoi22d1 U6068 ( .A1(n5821), .A2(n5803), .B1(n5802), .B2(n5804), .ZN(n5807)
         );
  aoi22d1 U6069 ( .A1(n5821), .A2(n5806), .B1(n5805), .B2(n5804), .ZN(n5842)
         );
  aoi22d1 U6070 ( .A1(n5862), .A2(n5807), .B1(n5842), .B2(n5830), .ZN(n5808)
         );
  oai22d1 U6071 ( .A1(n5877), .A2(n5809), .B1(n5910), .B2(n5808), .ZN(n5810)
         );
  aor211d1 U6072 ( .C1(n5881), .C2(n5812), .A(n5811), .B(n5810), .Z(n3157) );
  aoi22d1 U6073 ( .A1(n5885), .A2(mgmtsoc_litespisdrphycore_sr_out[25]), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[21]), .ZN(n5814) );
  aoi22d1 U6074 ( .A1(n5901), .A2(mgmtsoc_litespisdrphycore_sr_out[29]), .B1(
        n5886), .B2(mgmtsoc_litespisdrphycore_sr_out[27]), .ZN(n5813) );
  oai211d1 U6075 ( .C1(n5908), .C2(n5815), .A(n5814), .B(n5813), .ZN(n5826) );
  aoi22d1 U6076 ( .A1(n5821), .A2(n5817), .B1(n5816), .B2(n5818), .ZN(n5822)
         );
  aoi22d1 U6077 ( .A1(n5821), .A2(n5820), .B1(n5819), .B2(n5818), .ZN(n5851)
         );
  aoi22d1 U6078 ( .A1(n5862), .A2(n5822), .B1(n5851), .B2(n5830), .ZN(n5823)
         );
  oai22d1 U6079 ( .A1(n5877), .A2(n5824), .B1(n5910), .B2(n5823), .ZN(n5825)
         );
  aor211d1 U6080 ( .C1(n5881), .C2(n5827), .A(n5826), .B(n5825), .Z(n3156) );
  inv0d0 U6081 ( .I(mgmtsoc_litespisdrphycore_sr_out[26]), .ZN(n5840) );
  aoi22d1 U6082 ( .A1(n5893), .A2(mgmtsoc_litespisdrphycore_sr_out[23]), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[19]), .ZN(n5829) );
  aoi22d1 U6083 ( .A1(n5901), .A2(mgmtsoc_litespisdrphycore_sr_out[27]), .B1(
        n5886), .B2(mgmtsoc_litespisdrphycore_sr_out[25]), .ZN(n5828) );
  oai211d1 U6084 ( .C1(n5908), .C2(n5840), .A(n5829), .B(n5828), .ZN(n5836) );
  aoi22d1 U6085 ( .A1(n5862), .A2(n5832), .B1(n5831), .B2(n5830), .ZN(n5833)
         );
  oai22d1 U6086 ( .A1(n5877), .A2(n5834), .B1(n5910), .B2(n5833), .ZN(n5835)
         );
  aor211d1 U6087 ( .C1(n5881), .C2(n5837), .A(n5836), .B(n5835), .Z(n3154) );
  aoi22d1 U6088 ( .A1(n5893), .A2(mgmtsoc_litespisdrphycore_sr_out[22]), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[18]), .ZN(n5839) );
  aoi22d1 U6089 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[25]), .B1(
        n5886), .B2(mgmtsoc_litespisdrphycore_sr_out[24]), .ZN(n5838) );
  oai211d1 U6090 ( .C1(n5906), .C2(n5840), .A(n5839), .B(n5838), .ZN(n5846) );
  aoi22d1 U6091 ( .A1(n5862), .A2(n5842), .B1(n5841), .B2(n5863), .ZN(n5843)
         );
  oai22d1 U6092 ( .A1(n5877), .A2(n5844), .B1(n5910), .B2(n5843), .ZN(n5845)
         );
  aor211d1 U6093 ( .C1(n5881), .C2(n5847), .A(n5846), .B(n5845), .Z(n3153) );
  aoi22d1 U6094 ( .A1(n5893), .A2(mgmtsoc_litespisdrphycore_sr_out[21]), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[17]), .ZN(n5849) );
  aoi22d1 U6095 ( .A1(n5901), .A2(mgmtsoc_litespisdrphycore_sr_out[25]), .B1(
        n5897), .B2(mgmtsoc_litespisdrphycore_sr_out[23]), .ZN(n5848) );
  oai211d1 U6096 ( .C1(n5908), .C2(n5859), .A(n5849), .B(n5848), .ZN(n5855) );
  aoi22d1 U6097 ( .A1(n5862), .A2(n5851), .B1(n5850), .B2(n5863), .ZN(n5852)
         );
  oai22d1 U6098 ( .A1(n5877), .A2(n5853), .B1(n5910), .B2(n5852), .ZN(n5854)
         );
  aor211d1 U6099 ( .C1(n5881), .C2(n5856), .A(n5855), .B(n5854), .Z(n3152) );
  aoi22d1 U6100 ( .A1(n5897), .A2(mgmtsoc_litespisdrphycore_sr_out[22]), .B1(
        n5893), .B2(mgmtsoc_litespisdrphycore_sr_out[20]), .ZN(n5858) );
  aoi22d1 U6101 ( .A1(n5874), .A2(mgmtsoc_litespisdrphycore_sr_out[23]), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[16]), .ZN(n5857) );
  oai211d1 U6102 ( .C1(n5906), .C2(n5859), .A(n5858), .B(n5857), .ZN(n5868) );
  aoi22d1 U6103 ( .A1(n5862), .A2(n5861), .B1(n5860), .B2(n5863), .ZN(n5875)
         );
  aoi22d1 U6104 ( .A1(n5862), .A2(n5865), .B1(n5864), .B2(n5863), .ZN(n5866)
         );
  oai22d1 U6105 ( .A1(n5877), .A2(n5875), .B1(n5910), .B2(n5866), .ZN(n5867)
         );
  aor211d1 U6106 ( .C1(n5881), .C2(n5869), .A(n5868), .B(n5867), .Z(n3151) );
  aoi22d1 U6107 ( .A1(n5885), .A2(mgmtsoc_litespisdrphycore_sr_out[12]), .B1(
        n5870), .B2(mgmtsoc_litespisdrphycore_sr_out[8]), .ZN(n5873) );
  aoi22d1 U6108 ( .A1(n5871), .A2(mgmtsoc_litespisdrphycore_sr_out[16]), .B1(
        n5886), .B2(mgmtsoc_litespisdrphycore_sr_out[14]), .ZN(n5872) );
  oaim211d1 U6109 ( .C1(n5874), .C2(mgmtsoc_litespisdrphycore_sr_out[15]), .A(
        n5873), .B(n5872), .ZN(n5879) );
  oai22d1 U6110 ( .A1(n5877), .A2(n5876), .B1(n5910), .B2(n5875), .ZN(n5878)
         );
  aor211d1 U6111 ( .C1(n5881), .C2(n5880), .A(n5879), .B(n5878), .Z(n3143) );
  aoi22d1 U6112 ( .A1(n5897), .A2(mgmtsoc_litespisdrphycore_sr_out[5]), .B1(
        n5893), .B2(mgmtsoc_litespisdrphycore_sr_out[3]), .ZN(n5883) );
  aoi22d1 U6113 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[6]), .B1(
        n5901), .B2(mgmtsoc_litespisdrphycore_sr_out[7]), .ZN(n5882) );
  oai211d1 U6114 ( .C1(n5884), .C2(n5910), .A(n5883), .B(n5882), .ZN(n3134) );
  aoi22d1 U6115 ( .A1(n5886), .A2(mgmtsoc_litespisdrphycore_sr_out[4]), .B1(
        n5885), .B2(mgmtsoc_litespisdrphycore_sr_out[2]), .ZN(n5888) );
  aoi22d1 U6116 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[5]), .B1(
        n5901), .B2(mgmtsoc_litespisdrphycore_sr_out[6]), .ZN(n5887) );
  oai211d1 U6117 ( .C1(n5910), .C2(n5889), .A(n5888), .B(n5887), .ZN(n3133) );
  aoi22d1 U6118 ( .A1(n5897), .A2(mgmtsoc_litespisdrphycore_sr_out[3]), .B1(
        n5893), .B2(mgmtsoc_litespisdrphycore_sr_out[1]), .ZN(n5891) );
  aoi22d1 U6119 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[4]), .B1(
        n5901), .B2(mgmtsoc_litespisdrphycore_sr_out[5]), .ZN(n5890) );
  oai211d1 U6120 ( .C1(n5892), .C2(n5910), .A(n5891), .B(n5890), .ZN(n3132) );
  aoi22d1 U6121 ( .A1(n5897), .A2(mgmtsoc_litespisdrphycore_sr_out[2]), .B1(
        n5893), .B2(mgmtsoc_litespisdrphycore_sr_out[0]), .ZN(n5895) );
  aoi22d1 U6122 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[3]), .B1(
        n5901), .B2(mgmtsoc_litespisdrphycore_sr_out[4]), .ZN(n5894) );
  oai211d1 U6123 ( .C1(n5896), .C2(n5910), .A(n5895), .B(n5894), .ZN(n3131) );
  aoi22d1 U6124 ( .A1(n5901), .A2(mgmtsoc_litespisdrphycore_sr_out[3]), .B1(
        n5897), .B2(mgmtsoc_litespisdrphycore_sr_out[1]), .ZN(n5899) );
  nd02d0 U6125 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[2]), .ZN(
        n5898) );
  oai211d1 U6126 ( .C1(n5900), .C2(n5910), .A(n5899), .B(n5898), .ZN(n3130) );
  aoi22d1 U6127 ( .A1(n5902), .A2(mgmtsoc_litespisdrphycore_sr_out[1]), .B1(
        n5901), .B2(mgmtsoc_litespisdrphycore_sr_out[2]), .ZN(n5904) );
  nd02d0 U6128 ( .A1(n5886), .A2(mgmtsoc_litespisdrphycore_sr_out[0]), .ZN(
        n5903) );
  oai211d1 U6129 ( .C1(n5905), .C2(n5910), .A(n5904), .B(n5903), .ZN(n3129) );
  inv0d0 U6130 ( .I(mgmtsoc_litespisdrphycore_sr_out[1]), .ZN(n5907) );
  oai222d1 U6131 ( .A1(n5911), .A2(n5910), .B1(n5909), .B2(n5908), .C1(n5907), 
        .C2(n5906), .ZN(n3128) );
  nr13d1 U6132 ( .A1(n5915), .A2(n5914), .A3(n5926), .ZN(n5916) );
  mx02d1 U6133 ( .I0(n5917), .I1(mgmtsoc_litespisdrphycore_sr_cnt[1]), .S(
        n5916), .Z(n5918) );
  aoi22d1 U6134 ( .A1(n5941), .A2(n5919), .B1(n5918), .B2(n5951), .ZN(n3127)
         );
  nd03d0 U6135 ( .A1(n5925), .A2(mgmtsoc_litespisdrphycore_sr_cnt[0]), .A3(
        n5951), .ZN(n5924) );
  aon211d1 U6136 ( .C1(n5922), .C2(n5921), .B(n5920), .A(n5941), .ZN(n5923) );
  oai211d1 U6137 ( .C1(n5925), .C2(mgmtsoc_litespisdrphycore_sr_cnt[0]), .A(
        n5924), .B(n5923), .ZN(n3126) );
  aoi21d1 U6138 ( .B1(n5929), .B2(n5928), .A(n5926), .ZN(n5927) );
  oai21d1 U6139 ( .B1(n5929), .B2(n5928), .A(n5927), .ZN(n5935) );
  oai22d1 U6140 ( .A1(mgmtsoc_litespisdrphycore_sr_cnt[2]), .A2(n5935), .B1(
        n5951), .B2(n5933), .ZN(n5934) );
  aor31d1 U6141 ( .B1(n5951), .B2(mgmtsoc_litespisdrphycore_sr_cnt[2]), .B3(
        n5935), .A(n5934), .Z(n3125) );
  nd02d0 U6142 ( .A1(n5938), .A2(n5937), .ZN(n5936) );
  oai21d1 U6143 ( .B1(n5938), .B2(n5937), .A(n5936), .ZN(n5948) );
  oai21d1 U6144 ( .B1(n5949), .B2(n5948), .A(n5941), .ZN(n5947) );
  inv0d0 U6145 ( .I(n5939), .ZN(n5944) );
  oai22d1 U6146 ( .A1(n5942), .A2(n5945), .B1(n5941), .B2(n5940), .ZN(n5943)
         );
  oai21d1 U6147 ( .B1(n5945), .B2(n5944), .A(n5943), .ZN(n5946) );
  aon211d1 U6148 ( .C1(n5949), .C2(n5948), .B(n5947), .A(n5946), .ZN(n3124) );
  aoi31d1 U6149 ( .B1(mgmtsoc_litespisdrphycore_sr_cnt[7]), .B2(n5951), .B3(
        n5953), .A(n5950), .ZN(n5952) );
  oai21d1 U6150 ( .B1(mgmtsoc_litespisdrphycore_sr_cnt[7]), .B2(n5953), .A(
        n5952), .ZN(n3120) );
  inv0d0 U6151 ( .I(dbg_uart_cmd[0]), .ZN(n5958) );
  nd02d0 U6152 ( .A1(n5955), .A2(n5954), .ZN(n5966) );
  nd02d0 U6153 ( .A1(n5957), .A2(n5340), .ZN(n5965) );
  oai22d1 U6154 ( .A1(n5958), .A2(n5966), .B1(n5969), .B2(n5965), .ZN(n3117)
         );
  inv0d0 U6155 ( .I(dbg_uart_cmd[1]), .ZN(n5959) );
  oai22d1 U6156 ( .A1(n5959), .A2(n5966), .B1(n5970), .B2(n5965), .ZN(n3116)
         );
  oai22d1 U6157 ( .A1(n5960), .A2(n5966), .B1(n5971), .B2(n5965), .ZN(n3115)
         );
  inv0d0 U6158 ( .I(dbg_uart_cmd[3]), .ZN(n5961) );
  oai22d1 U6159 ( .A1(n5961), .A2(n5966), .B1(n5972), .B2(n5965), .ZN(n3114)
         );
  inv0d0 U6160 ( .I(dbg_uart_cmd[4]), .ZN(n5962) );
  oai22d1 U6161 ( .A1(n5962), .A2(n5966), .B1(n5973), .B2(n5965), .ZN(n3113)
         );
  inv0d0 U6162 ( .I(dbg_uart_cmd[5]), .ZN(n5963) );
  oai22d1 U6163 ( .A1(n5963), .A2(n5966), .B1(n5974), .B2(n5965), .ZN(n3112)
         );
  oai22d1 U6164 ( .A1(n5964), .A2(n5966), .B1(n5975), .B2(n5965), .ZN(n3111)
         );
  oai22d1 U6165 ( .A1(n5967), .A2(n5966), .B1(n5976), .B2(n5965), .ZN(n3110)
         );
  inv0d1 U6166 ( .I(n5968), .ZN(n5977) );
  aoim22d1 U6167 ( .A1(n5977), .A2(n5969), .B1(dbg_uart_length[0]), .B2(n5977), 
        .Z(n3109) );
  aoim22d1 U6168 ( .A1(n5977), .A2(n5970), .B1(dbg_uart_length[1]), .B2(n5977), 
        .Z(n3108) );
  aoim22d1 U6169 ( .A1(n5977), .A2(n5971), .B1(dbg_uart_length[2]), .B2(n5977), 
        .Z(n3107) );
  aoim22d1 U6170 ( .A1(n5977), .A2(n5972), .B1(dbg_uart_length[3]), .B2(n5977), 
        .Z(n3106) );
  aoim22d1 U6171 ( .A1(n5977), .A2(n5973), .B1(dbg_uart_length[4]), .B2(n5977), 
        .Z(n3105) );
  aoim22d1 U6172 ( .A1(n5977), .A2(n5974), .B1(dbg_uart_length[5]), .B2(n5977), 
        .Z(n3104) );
  aoim22d1 U6173 ( .A1(n5977), .A2(n5975), .B1(dbg_uart_length[6]), .B2(n5977), 
        .Z(n3103) );
  aoim22d1 U6174 ( .A1(n5977), .A2(n5976), .B1(dbg_uart_length[7]), .B2(n5977), 
        .Z(n3102) );
  inv0d0 U6175 ( .I(n5979), .ZN(n5980) );
  aoim211d1 U6176 ( .C1(dbg_uart_tx_tick), .C2(dbg_uart_tx_count[0]), .A(n5980), .B(n5990), .ZN(n3101) );
  inv0d0 U6177 ( .I(dbg_uart_tx_count[1]), .ZN(n5978) );
  nr02d0 U6178 ( .A1(n5979), .A2(n5978), .ZN(n5981) );
  aoi211d1 U6179 ( .C1(n5979), .C2(n5978), .A(n5981), .B(n5990), .ZN(n3100) );
  nd03d0 U6180 ( .A1(n5980), .A2(dbg_uart_tx_count[2]), .A3(
        dbg_uart_tx_count[1]), .ZN(n5983) );
  ora211d1 U6181 ( .C1(dbg_uart_tx_count[2]), .C2(n5981), .A(n5983), .B(n5987), 
        .Z(n3099) );
  nr02d0 U6182 ( .A1(n5984), .A2(n5983), .ZN(n5982) );
  aoi211d1 U6183 ( .C1(n5984), .C2(n5983), .A(n5990), .B(n5982), .ZN(n3098) );
  oai21d1 U6184 ( .B1(n5985), .B2(n5990), .A(n6019), .ZN(n3097) );
  inv0d0 U6185 ( .I(n5986), .ZN(n6015) );
  aoi22d1 U6186 ( .A1(dbg_uart_wishbone_dat_w[0]), .A2(n6015), .B1(
        dbg_uart_wishbone_dat_w[8]), .B2(n6013), .ZN(n5993) );
  nr02d0 U6187 ( .A1(dbg_uart_bytes_count[0]), .A2(dbg_uart_bytes_count[1]), 
        .ZN(n6014) );
  aoi22d1 U6188 ( .A1(dbg_uart_wishbone_dat_w[16]), .A2(n6012), .B1(
        dbg_uart_wishbone_dat_w[24]), .B2(n6014), .ZN(n5992) );
  an02d0 U6189 ( .A1(dbg_uart_tx_tick), .A2(n5987), .Z(n6016) );
  oai22d1 U6190 ( .A1(dbg_uart_tx_tick), .A2(n5990), .B1(n5989), .B2(n5988), 
        .ZN(n6017) );
  aoi22d1 U6191 ( .A1(dbg_uart_tx_data[1]), .A2(n6016), .B1(
        dbg_uart_tx_data[0]), .B2(n6017), .ZN(n5991) );
  aon211d1 U6192 ( .C1(n5993), .C2(n5992), .B(n6019), .A(n5991), .ZN(n3096) );
  aoi22d1 U6193 ( .A1(dbg_uart_wishbone_dat_w[1]), .A2(n6015), .B1(
        dbg_uart_wishbone_dat_w[25]), .B2(n6014), .ZN(n5996) );
  aoi22d1 U6194 ( .A1(dbg_uart_wishbone_dat_w[9]), .A2(n6013), .B1(
        dbg_uart_wishbone_dat_w[17]), .B2(n6012), .ZN(n5995) );
  aoi22d1 U6195 ( .A1(dbg_uart_tx_data[2]), .A2(n6016), .B1(
        dbg_uart_tx_data[1]), .B2(n6017), .ZN(n5994) );
  aon211d1 U6196 ( .C1(n5996), .C2(n5995), .B(n6019), .A(n5994), .ZN(n3095) );
  aoi22d1 U6197 ( .A1(dbg_uart_wishbone_dat_w[2]), .A2(n6015), .B1(
        dbg_uart_wishbone_dat_w[26]), .B2(n6014), .ZN(n5999) );
  aoi22d1 U6198 ( .A1(dbg_uart_wishbone_dat_w[10]), .A2(n6013), .B1(
        dbg_uart_wishbone_dat_w[18]), .B2(n6012), .ZN(n5998) );
  aoi22d1 U6199 ( .A1(dbg_uart_tx_data[3]), .A2(n6016), .B1(
        dbg_uart_tx_data[2]), .B2(n6017), .ZN(n5997) );
  aon211d1 U6200 ( .C1(n5999), .C2(n5998), .B(n6019), .A(n5997), .ZN(n3094) );
  aoi22d1 U6201 ( .A1(dbg_uart_wishbone_dat_w[3]), .A2(n6015), .B1(
        dbg_uart_wishbone_dat_w[19]), .B2(n6012), .ZN(n6002) );
  aoi22d1 U6202 ( .A1(dbg_uart_wishbone_dat_w[11]), .A2(n6013), .B1(
        dbg_uart_wishbone_dat_w[27]), .B2(n6014), .ZN(n6001) );
  aoi22d1 U6203 ( .A1(dbg_uart_tx_data[4]), .A2(n6016), .B1(
        dbg_uart_tx_data[3]), .B2(n6017), .ZN(n6000) );
  aon211d1 U6204 ( .C1(n6002), .C2(n6001), .B(n6019), .A(n6000), .ZN(n3093) );
  aoi22d1 U6205 ( .A1(dbg_uart_wishbone_dat_w[20]), .A2(n6012), .B1(
        dbg_uart_wishbone_dat_w[28]), .B2(n6014), .ZN(n6005) );
  aoi22d1 U6206 ( .A1(dbg_uart_wishbone_dat_w[4]), .A2(n6015), .B1(
        dbg_uart_wishbone_dat_w[12]), .B2(n6013), .ZN(n6004) );
  aoi22d1 U6207 ( .A1(dbg_uart_tx_data[5]), .A2(n6016), .B1(
        dbg_uart_tx_data[4]), .B2(n6017), .ZN(n6003) );
  aon211d1 U6208 ( .C1(n6005), .C2(n6004), .B(n6019), .A(n6003), .ZN(n3092) );
  aoi22d1 U6209 ( .A1(dbg_uart_wishbone_dat_w[13]), .A2(n6013), .B1(
        dbg_uart_wishbone_dat_w[29]), .B2(n6014), .ZN(n6008) );
  aoi22d1 U6210 ( .A1(dbg_uart_wishbone_dat_w[5]), .A2(n6015), .B1(
        dbg_uart_wishbone_dat_w[21]), .B2(n6012), .ZN(n6007) );
  aoi22d1 U6211 ( .A1(dbg_uart_tx_data[6]), .A2(n6016), .B1(
        dbg_uart_tx_data[5]), .B2(n6017), .ZN(n6006) );
  aon211d1 U6212 ( .C1(n6008), .C2(n6007), .B(n6019), .A(n6006), .ZN(n3091) );
  aoi22d1 U6213 ( .A1(dbg_uart_wishbone_dat_w[6]), .A2(n6015), .B1(
        dbg_uart_wishbone_dat_w[14]), .B2(n6013), .ZN(n6011) );
  aoi22d1 U6214 ( .A1(dbg_uart_wishbone_dat_w[22]), .A2(n6012), .B1(
        dbg_uart_wishbone_dat_w[30]), .B2(n6014), .ZN(n6010) );
  aoi22d1 U6215 ( .A1(dbg_uart_tx_data[7]), .A2(n6016), .B1(
        dbg_uart_tx_data[6]), .B2(n6017), .ZN(n6009) );
  aon211d1 U6216 ( .C1(n6011), .C2(n6010), .B(n6019), .A(n6009), .ZN(n3090) );
  aoi22d1 U6217 ( .A1(dbg_uart_wishbone_dat_w[15]), .A2(n6013), .B1(
        dbg_uart_wishbone_dat_w[23]), .B2(n6012), .ZN(n6021) );
  aoi22d1 U6218 ( .A1(dbg_uart_wishbone_dat_w[7]), .A2(n6015), .B1(
        dbg_uart_wishbone_dat_w[31]), .B2(n6014), .ZN(n6020) );
  aoi21d1 U6219 ( .B1(dbg_uart_tx_data[7]), .B2(n6017), .A(n6016), .ZN(n6018)
         );
  aon211d1 U6220 ( .C1(n6021), .C2(n6020), .B(n6019), .A(n6018), .ZN(n3088) );
endmodule

