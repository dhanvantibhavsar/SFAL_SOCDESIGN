module VexRiscv ( vccd1, vssd1, externalResetVector, timerInterrupt, 
        softwareInterrupt, externalInterruptArray, debug_bus_cmd_valid, 
        debug_bus_cmd_ready, debug_bus_cmd_payload_wr, 
        debug_bus_cmd_payload_address, debug_bus_cmd_payload_data, 
        debug_bus_rsp_data, debug_resetOut, iBusWishbone_CYC, iBusWishbone_STB, 
        iBusWishbone_ACK, iBusWishbone_WE, iBusWishbone_DAT_MISO, 
        iBusWishbone_DAT_MOSI, iBusWishbone_SEL, iBusWishbone_ERR, 
        iBusWishbone_CTI, iBusWishbone_BTE, dBusWishbone_CYC, dBusWishbone_STB, 
        dBusWishbone_ACK, dBusWishbone_WE, dBusWishbone_ADR, 
        dBusWishbone_DAT_MISO, dBusWishbone_DAT_MOSI, dBusWishbone_SEL, 
        dBusWishbone_ERR, dBusWishbone_CTI, dBusWishbone_BTE, clk, reset, 
        debugReset, \iBusWishbone_ADR[29] , \iBusWishbone_ADR[28] , 
        \iBusWishbone_ADR[27] , \iBusWishbone_ADR[26] , \iBusWishbone_ADR[25] , 
        \iBusWishbone_ADR[24] , \iBusWishbone_ADR[23] , \iBusWishbone_ADR[22] , 
        \iBusWishbone_ADR[21] , \iBusWishbone_ADR[20] , \iBusWishbone_ADR[19] , 
        \iBusWishbone_ADR[18] , \iBusWishbone_ADR[17] , \iBusWishbone_ADR[16] , 
        \iBusWishbone_ADR[15] , \iBusWishbone_ADR[14] , \iBusWishbone_ADR[13] , 
        \iBusWishbone_ADR[12] , \iBusWishbone_ADR[11] , \iBusWishbone_ADR[10] , 
        \iBusWishbone_ADR[9] , \iBusWishbone_ADR[8] , \iBusWishbone_ADR[7] , 
        \iBusWishbone_ADR[6] , \iBusWishbone_ADR[5] , \iBusWishbone_ADR[4] , 
        \iBusWishbone_ADR[3]_BAR , \iBusWishbone_ADR[2] , 
        \iBusWishbone_ADR[1] , \iBusWishbone_ADR[0]  );
  input [31:0] externalResetVector;
  input [31:0] externalInterruptArray;
  input [7:0] debug_bus_cmd_payload_address;
  input [31:0] debug_bus_cmd_payload_data;
  output [31:0] debug_bus_rsp_data;
  input [31:0] iBusWishbone_DAT_MISO;
  output [31:0] iBusWishbone_DAT_MOSI;
  output [3:0] iBusWishbone_SEL;
  output [2:0] iBusWishbone_CTI;
  output [1:0] iBusWishbone_BTE;
  output [29:0] dBusWishbone_ADR;
  input [31:0] dBusWishbone_DAT_MISO;
  output [31:0] dBusWishbone_DAT_MOSI;
  output [3:0] dBusWishbone_SEL;
  output [2:0] dBusWishbone_CTI;
  output [1:0] dBusWishbone_BTE;
  input timerInterrupt, softwareInterrupt, debug_bus_cmd_valid,
         debug_bus_cmd_payload_wr, iBusWishbone_ACK, iBusWishbone_ERR,
         dBusWishbone_ACK, dBusWishbone_ERR, clk, reset, debugReset;
  output debug_bus_cmd_ready, debug_resetOut, iBusWishbone_CYC,
         iBusWishbone_STB, iBusWishbone_WE, dBusWishbone_CYC, dBusWishbone_STB,
         dBusWishbone_WE, \iBusWishbone_ADR[29] , \iBusWishbone_ADR[28] ,
         \iBusWishbone_ADR[27] , \iBusWishbone_ADR[26] ,
         \iBusWishbone_ADR[25] , \iBusWishbone_ADR[24] ,
         \iBusWishbone_ADR[23] , \iBusWishbone_ADR[22] ,
         \iBusWishbone_ADR[21] , \iBusWishbone_ADR[20] ,
         \iBusWishbone_ADR[19] , \iBusWishbone_ADR[18] ,
         \iBusWishbone_ADR[17] , \iBusWishbone_ADR[16] ,
         \iBusWishbone_ADR[15] , \iBusWishbone_ADR[14] ,
         \iBusWishbone_ADR[13] , \iBusWishbone_ADR[12] ,
         \iBusWishbone_ADR[11] , \iBusWishbone_ADR[10] , \iBusWishbone_ADR[9] ,
         \iBusWishbone_ADR[8] , \iBusWishbone_ADR[7] , \iBusWishbone_ADR[6] ,
         \iBusWishbone_ADR[5] , \iBusWishbone_ADR[4] ,
         \iBusWishbone_ADR[3]_BAR , \iBusWishbone_ADR[2] ,
         \iBusWishbone_ADR[1] , \iBusWishbone_ADR[0] ;
  inout vccd1,  vssd1;
  wire   n7265, \_zz_IBusCachedPlugin_fetchPc_pc_1[2] , memory_MEMORY_STORE,
         execute_SRC_USE_SUB_LESS, _zz__zz_execute_BranchPlugin_branch_src2_3,
         _zz__zz_execute_BranchPlugin_branch_src2_2,
         _zz__zz_execute_BranchPlugin_branch_src2_1,
         _zz__zz_execute_BranchPlugin_branch_src2_0, decode_INSTRUCTION_30,
         decode_INSTRUCTION_24, decode_INSTRUCTION_23, decode_INSTRUCTION_22,
         decode_INSTRUCTION_21, decode_INSTRUCTION_11, decode_INSTRUCTION_10,
         decode_INSTRUCTION_9, decode_INSTRUCTION_8, decode_INSTRUCTION_7,
         _zz_decode_LEGAL_INSTRUCTION_1_13,
         \_zz_decode_LEGAL_INSTRUCTION_7[14] ,
         _zz_decode_LEGAL_INSTRUCTION_7_12, _zz_decode_LEGAL_INSTRUCTION_13_31,
         \_zz__zz_decode_ENV_CTRL_2_1[20] , \RegFilePlugin_regFile[0][31] ,
         \RegFilePlugin_regFile[0][30] , \RegFilePlugin_regFile[0][29] ,
         \RegFilePlugin_regFile[0][28] , \RegFilePlugin_regFile[0][27] ,
         \RegFilePlugin_regFile[0][26] , \RegFilePlugin_regFile[0][25] ,
         \RegFilePlugin_regFile[0][24] , \RegFilePlugin_regFile[0][23] ,
         \RegFilePlugin_regFile[0][22] , \RegFilePlugin_regFile[0][21] ,
         \RegFilePlugin_regFile[0][20] , \RegFilePlugin_regFile[0][19] ,
         \RegFilePlugin_regFile[0][18] , \RegFilePlugin_regFile[0][17] ,
         \RegFilePlugin_regFile[0][16] , \RegFilePlugin_regFile[0][15] ,
         \RegFilePlugin_regFile[0][14] , \RegFilePlugin_regFile[0][13] ,
         \RegFilePlugin_regFile[0][12] , \RegFilePlugin_regFile[0][11] ,
         \RegFilePlugin_regFile[0][10] , \RegFilePlugin_regFile[0][9] ,
         \RegFilePlugin_regFile[0][8] , \RegFilePlugin_regFile[0][7] ,
         \RegFilePlugin_regFile[0][6] , \RegFilePlugin_regFile[0][5] ,
         \RegFilePlugin_regFile[0][4] , \RegFilePlugin_regFile[0][3] ,
         \RegFilePlugin_regFile[0][2] , \RegFilePlugin_regFile[0][1] ,
         \RegFilePlugin_regFile[0][0] , \RegFilePlugin_regFile[1][31] ,
         \RegFilePlugin_regFile[1][30] , \RegFilePlugin_regFile[1][29] ,
         \RegFilePlugin_regFile[1][28] , \RegFilePlugin_regFile[1][27] ,
         \RegFilePlugin_regFile[1][26] , \RegFilePlugin_regFile[1][25] ,
         \RegFilePlugin_regFile[1][24] , \RegFilePlugin_regFile[1][23] ,
         \RegFilePlugin_regFile[1][22] , \RegFilePlugin_regFile[1][21] ,
         \RegFilePlugin_regFile[1][20] , \RegFilePlugin_regFile[1][19] ,
         \RegFilePlugin_regFile[1][18] , \RegFilePlugin_regFile[1][17] ,
         \RegFilePlugin_regFile[1][16] , \RegFilePlugin_regFile[1][15] ,
         \RegFilePlugin_regFile[1][14] , \RegFilePlugin_regFile[1][13] ,
         \RegFilePlugin_regFile[1][12] , \RegFilePlugin_regFile[1][11] ,
         \RegFilePlugin_regFile[1][10] , \RegFilePlugin_regFile[1][9] ,
         \RegFilePlugin_regFile[1][8] , \RegFilePlugin_regFile[1][7] ,
         \RegFilePlugin_regFile[1][6] , \RegFilePlugin_regFile[1][5] ,
         \RegFilePlugin_regFile[1][4] , \RegFilePlugin_regFile[1][3] ,
         \RegFilePlugin_regFile[1][2] , \RegFilePlugin_regFile[1][1] ,
         \RegFilePlugin_regFile[1][0] , \RegFilePlugin_regFile[2][31] ,
         \RegFilePlugin_regFile[2][30] , \RegFilePlugin_regFile[2][29] ,
         \RegFilePlugin_regFile[2][28] , \RegFilePlugin_regFile[2][27] ,
         \RegFilePlugin_regFile[2][26] , \RegFilePlugin_regFile[2][25] ,
         \RegFilePlugin_regFile[2][24] , \RegFilePlugin_regFile[2][23] ,
         \RegFilePlugin_regFile[2][22] , \RegFilePlugin_regFile[2][21] ,
         \RegFilePlugin_regFile[2][20] , \RegFilePlugin_regFile[2][19] ,
         \RegFilePlugin_regFile[2][18] , \RegFilePlugin_regFile[2][17] ,
         \RegFilePlugin_regFile[2][16] , \RegFilePlugin_regFile[2][15] ,
         \RegFilePlugin_regFile[2][14] , \RegFilePlugin_regFile[2][13] ,
         \RegFilePlugin_regFile[2][12] , \RegFilePlugin_regFile[2][11] ,
         \RegFilePlugin_regFile[2][10] , \RegFilePlugin_regFile[2][9] ,
         \RegFilePlugin_regFile[2][8] , \RegFilePlugin_regFile[2][7] ,
         \RegFilePlugin_regFile[2][6] , \RegFilePlugin_regFile[2][5] ,
         \RegFilePlugin_regFile[2][4] , \RegFilePlugin_regFile[2][3] ,
         \RegFilePlugin_regFile[2][2] , \RegFilePlugin_regFile[2][1] ,
         \RegFilePlugin_regFile[2][0] , \RegFilePlugin_regFile[3][31] ,
         \RegFilePlugin_regFile[3][30] , \RegFilePlugin_regFile[3][29] ,
         \RegFilePlugin_regFile[3][28] , \RegFilePlugin_regFile[3][27] ,
         \RegFilePlugin_regFile[3][26] , \RegFilePlugin_regFile[3][25] ,
         \RegFilePlugin_regFile[3][24] , \RegFilePlugin_regFile[3][23] ,
         \RegFilePlugin_regFile[3][22] , \RegFilePlugin_regFile[3][21] ,
         \RegFilePlugin_regFile[3][20] , \RegFilePlugin_regFile[3][19] ,
         \RegFilePlugin_regFile[3][18] , \RegFilePlugin_regFile[3][17] ,
         \RegFilePlugin_regFile[3][16] , \RegFilePlugin_regFile[3][15] ,
         \RegFilePlugin_regFile[3][14] , \RegFilePlugin_regFile[3][13] ,
         \RegFilePlugin_regFile[3][12] , \RegFilePlugin_regFile[3][11] ,
         \RegFilePlugin_regFile[3][10] , \RegFilePlugin_regFile[3][9] ,
         \RegFilePlugin_regFile[3][8] , \RegFilePlugin_regFile[3][7] ,
         \RegFilePlugin_regFile[3][6] , \RegFilePlugin_regFile[3][5] ,
         \RegFilePlugin_regFile[3][4] , \RegFilePlugin_regFile[3][3] ,
         \RegFilePlugin_regFile[3][2] , \RegFilePlugin_regFile[3][1] ,
         \RegFilePlugin_regFile[3][0] , \RegFilePlugin_regFile[4][31] ,
         \RegFilePlugin_regFile[4][30] , \RegFilePlugin_regFile[4][29] ,
         \RegFilePlugin_regFile[4][28] , \RegFilePlugin_regFile[4][27] ,
         \RegFilePlugin_regFile[4][26] , \RegFilePlugin_regFile[4][25] ,
         \RegFilePlugin_regFile[4][24] , \RegFilePlugin_regFile[4][23] ,
         \RegFilePlugin_regFile[4][22] , \RegFilePlugin_regFile[4][21] ,
         \RegFilePlugin_regFile[4][20] , \RegFilePlugin_regFile[4][19] ,
         \RegFilePlugin_regFile[4][18] , \RegFilePlugin_regFile[4][17] ,
         \RegFilePlugin_regFile[4][16] , \RegFilePlugin_regFile[4][15] ,
         \RegFilePlugin_regFile[4][14] , \RegFilePlugin_regFile[4][13] ,
         \RegFilePlugin_regFile[4][12] , \RegFilePlugin_regFile[4][11] ,
         \RegFilePlugin_regFile[4][10] , \RegFilePlugin_regFile[4][9] ,
         \RegFilePlugin_regFile[4][8] , \RegFilePlugin_regFile[4][7] ,
         \RegFilePlugin_regFile[4][6] , \RegFilePlugin_regFile[4][5] ,
         \RegFilePlugin_regFile[4][4] , \RegFilePlugin_regFile[4][3] ,
         \RegFilePlugin_regFile[4][2] , \RegFilePlugin_regFile[4][1] ,
         \RegFilePlugin_regFile[4][0] , \RegFilePlugin_regFile[5][31] ,
         \RegFilePlugin_regFile[5][30] , \RegFilePlugin_regFile[5][29] ,
         \RegFilePlugin_regFile[5][28] , \RegFilePlugin_regFile[5][27] ,
         \RegFilePlugin_regFile[5][26] , \RegFilePlugin_regFile[5][25] ,
         \RegFilePlugin_regFile[5][24] , \RegFilePlugin_regFile[5][23] ,
         \RegFilePlugin_regFile[5][22] , \RegFilePlugin_regFile[5][21] ,
         \RegFilePlugin_regFile[5][20] , \RegFilePlugin_regFile[5][19] ,
         \RegFilePlugin_regFile[5][18] , \RegFilePlugin_regFile[5][17] ,
         \RegFilePlugin_regFile[5][16] , \RegFilePlugin_regFile[5][15] ,
         \RegFilePlugin_regFile[5][14] , \RegFilePlugin_regFile[5][13] ,
         \RegFilePlugin_regFile[5][12] , \RegFilePlugin_regFile[5][11] ,
         \RegFilePlugin_regFile[5][10] , \RegFilePlugin_regFile[5][9] ,
         \RegFilePlugin_regFile[5][8] , \RegFilePlugin_regFile[5][7] ,
         \RegFilePlugin_regFile[5][6] , \RegFilePlugin_regFile[5][5] ,
         \RegFilePlugin_regFile[5][4] , \RegFilePlugin_regFile[5][3] ,
         \RegFilePlugin_regFile[5][2] , \RegFilePlugin_regFile[5][1] ,
         \RegFilePlugin_regFile[5][0] , \RegFilePlugin_regFile[6][31] ,
         \RegFilePlugin_regFile[6][30] , \RegFilePlugin_regFile[6][29] ,
         \RegFilePlugin_regFile[6][28] , \RegFilePlugin_regFile[6][27] ,
         \RegFilePlugin_regFile[6][26] , \RegFilePlugin_regFile[6][25] ,
         \RegFilePlugin_regFile[6][24] , \RegFilePlugin_regFile[6][23] ,
         \RegFilePlugin_regFile[6][22] , \RegFilePlugin_regFile[6][21] ,
         \RegFilePlugin_regFile[6][20] , \RegFilePlugin_regFile[6][19] ,
         \RegFilePlugin_regFile[6][18] , \RegFilePlugin_regFile[6][17] ,
         \RegFilePlugin_regFile[6][16] , \RegFilePlugin_regFile[6][15] ,
         \RegFilePlugin_regFile[6][14] , \RegFilePlugin_regFile[6][13] ,
         \RegFilePlugin_regFile[6][12] , \RegFilePlugin_regFile[6][11] ,
         \RegFilePlugin_regFile[6][10] , \RegFilePlugin_regFile[6][9] ,
         \RegFilePlugin_regFile[6][8] , \RegFilePlugin_regFile[6][7] ,
         \RegFilePlugin_regFile[6][6] , \RegFilePlugin_regFile[6][5] ,
         \RegFilePlugin_regFile[6][4] , \RegFilePlugin_regFile[6][3] ,
         \RegFilePlugin_regFile[6][2] , \RegFilePlugin_regFile[6][1] ,
         \RegFilePlugin_regFile[6][0] , \RegFilePlugin_regFile[7][31] ,
         \RegFilePlugin_regFile[7][30] , \RegFilePlugin_regFile[7][29] ,
         \RegFilePlugin_regFile[7][28] , \RegFilePlugin_regFile[7][27] ,
         \RegFilePlugin_regFile[7][26] , \RegFilePlugin_regFile[7][25] ,
         \RegFilePlugin_regFile[7][24] , \RegFilePlugin_regFile[7][23] ,
         \RegFilePlugin_regFile[7][22] , \RegFilePlugin_regFile[7][21] ,
         \RegFilePlugin_regFile[7][20] , \RegFilePlugin_regFile[7][19] ,
         \RegFilePlugin_regFile[7][18] , \RegFilePlugin_regFile[7][17] ,
         \RegFilePlugin_regFile[7][16] , \RegFilePlugin_regFile[7][15] ,
         \RegFilePlugin_regFile[7][14] , \RegFilePlugin_regFile[7][13] ,
         \RegFilePlugin_regFile[7][12] , \RegFilePlugin_regFile[7][11] ,
         \RegFilePlugin_regFile[7][10] , \RegFilePlugin_regFile[7][9] ,
         \RegFilePlugin_regFile[7][8] , \RegFilePlugin_regFile[7][7] ,
         \RegFilePlugin_regFile[7][6] , \RegFilePlugin_regFile[7][5] ,
         \RegFilePlugin_regFile[7][4] , \RegFilePlugin_regFile[7][3] ,
         \RegFilePlugin_regFile[7][2] , \RegFilePlugin_regFile[7][1] ,
         \RegFilePlugin_regFile[7][0] , \RegFilePlugin_regFile[8][31] ,
         \RegFilePlugin_regFile[8][30] , \RegFilePlugin_regFile[8][29] ,
         \RegFilePlugin_regFile[8][28] , \RegFilePlugin_regFile[8][27] ,
         \RegFilePlugin_regFile[8][26] , \RegFilePlugin_regFile[8][25] ,
         \RegFilePlugin_regFile[8][24] , \RegFilePlugin_regFile[8][23] ,
         \RegFilePlugin_regFile[8][22] , \RegFilePlugin_regFile[8][21] ,
         \RegFilePlugin_regFile[8][20] , \RegFilePlugin_regFile[8][19] ,
         \RegFilePlugin_regFile[8][18] , \RegFilePlugin_regFile[8][17] ,
         \RegFilePlugin_regFile[8][16] , \RegFilePlugin_regFile[8][15] ,
         \RegFilePlugin_regFile[8][14] , \RegFilePlugin_regFile[8][13] ,
         \RegFilePlugin_regFile[8][12] , \RegFilePlugin_regFile[8][11] ,
         \RegFilePlugin_regFile[8][10] , \RegFilePlugin_regFile[8][9] ,
         \RegFilePlugin_regFile[8][8] , \RegFilePlugin_regFile[8][7] ,
         \RegFilePlugin_regFile[8][6] , \RegFilePlugin_regFile[8][5] ,
         \RegFilePlugin_regFile[8][4] , \RegFilePlugin_regFile[8][3] ,
         \RegFilePlugin_regFile[8][2] , \RegFilePlugin_regFile[8][1] ,
         \RegFilePlugin_regFile[8][0] , \RegFilePlugin_regFile[9][31] ,
         \RegFilePlugin_regFile[9][30] , \RegFilePlugin_regFile[9][29] ,
         \RegFilePlugin_regFile[9][28] , \RegFilePlugin_regFile[9][27] ,
         \RegFilePlugin_regFile[9][26] , \RegFilePlugin_regFile[9][25] ,
         \RegFilePlugin_regFile[9][24] , \RegFilePlugin_regFile[9][23] ,
         \RegFilePlugin_regFile[9][22] , \RegFilePlugin_regFile[9][21] ,
         \RegFilePlugin_regFile[9][20] , \RegFilePlugin_regFile[9][19] ,
         \RegFilePlugin_regFile[9][18] , \RegFilePlugin_regFile[9][17] ,
         \RegFilePlugin_regFile[9][16] , \RegFilePlugin_regFile[9][15] ,
         \RegFilePlugin_regFile[9][14] , \RegFilePlugin_regFile[9][13] ,
         \RegFilePlugin_regFile[9][12] , \RegFilePlugin_regFile[9][11] ,
         \RegFilePlugin_regFile[9][10] , \RegFilePlugin_regFile[9][9] ,
         \RegFilePlugin_regFile[9][8] , \RegFilePlugin_regFile[9][7] ,
         \RegFilePlugin_regFile[9][6] , \RegFilePlugin_regFile[9][5] ,
         \RegFilePlugin_regFile[9][4] , \RegFilePlugin_regFile[9][3] ,
         \RegFilePlugin_regFile[9][2] , \RegFilePlugin_regFile[9][1] ,
         \RegFilePlugin_regFile[9][0] , \RegFilePlugin_regFile[10][31] ,
         \RegFilePlugin_regFile[10][30] , \RegFilePlugin_regFile[10][29] ,
         \RegFilePlugin_regFile[10][28] , \RegFilePlugin_regFile[10][27] ,
         \RegFilePlugin_regFile[10][26] , \RegFilePlugin_regFile[10][25] ,
         \RegFilePlugin_regFile[10][24] , \RegFilePlugin_regFile[10][23] ,
         \RegFilePlugin_regFile[10][22] , \RegFilePlugin_regFile[10][21] ,
         \RegFilePlugin_regFile[10][20] , \RegFilePlugin_regFile[10][19] ,
         \RegFilePlugin_regFile[10][18] , \RegFilePlugin_regFile[10][17] ,
         \RegFilePlugin_regFile[10][16] , \RegFilePlugin_regFile[10][15] ,
         \RegFilePlugin_regFile[10][14] , \RegFilePlugin_regFile[10][13] ,
         \RegFilePlugin_regFile[10][12] , \RegFilePlugin_regFile[10][11] ,
         \RegFilePlugin_regFile[10][10] , \RegFilePlugin_regFile[10][9] ,
         \RegFilePlugin_regFile[10][8] , \RegFilePlugin_regFile[10][7] ,
         \RegFilePlugin_regFile[10][6] , \RegFilePlugin_regFile[10][5] ,
         \RegFilePlugin_regFile[10][4] , \RegFilePlugin_regFile[10][3] ,
         \RegFilePlugin_regFile[10][2] , \RegFilePlugin_regFile[10][1] ,
         \RegFilePlugin_regFile[10][0] , \RegFilePlugin_regFile[11][31] ,
         \RegFilePlugin_regFile[11][30] , \RegFilePlugin_regFile[11][29] ,
         \RegFilePlugin_regFile[11][28] , \RegFilePlugin_regFile[11][27] ,
         \RegFilePlugin_regFile[11][26] , \RegFilePlugin_regFile[11][25] ,
         \RegFilePlugin_regFile[11][24] , \RegFilePlugin_regFile[11][23] ,
         \RegFilePlugin_regFile[11][22] , \RegFilePlugin_regFile[11][21] ,
         \RegFilePlugin_regFile[11][20] , \RegFilePlugin_regFile[11][19] ,
         \RegFilePlugin_regFile[11][18] , \RegFilePlugin_regFile[11][17] ,
         \RegFilePlugin_regFile[11][16] , \RegFilePlugin_regFile[11][15] ,
         \RegFilePlugin_regFile[11][14] , \RegFilePlugin_regFile[11][13] ,
         \RegFilePlugin_regFile[11][12] , \RegFilePlugin_regFile[11][11] ,
         \RegFilePlugin_regFile[11][10] , \RegFilePlugin_regFile[11][9] ,
         \RegFilePlugin_regFile[11][8] , \RegFilePlugin_regFile[11][7] ,
         \RegFilePlugin_regFile[11][6] , \RegFilePlugin_regFile[11][5] ,
         \RegFilePlugin_regFile[11][4] , \RegFilePlugin_regFile[11][3] ,
         \RegFilePlugin_regFile[11][2] , \RegFilePlugin_regFile[11][1] ,
         \RegFilePlugin_regFile[11][0] , \RegFilePlugin_regFile[12][31] ,
         \RegFilePlugin_regFile[12][30] , \RegFilePlugin_regFile[12][29] ,
         \RegFilePlugin_regFile[12][28] , \RegFilePlugin_regFile[12][27] ,
         \RegFilePlugin_regFile[12][26] , \RegFilePlugin_regFile[12][25] ,
         \RegFilePlugin_regFile[12][24] , \RegFilePlugin_regFile[12][23] ,
         \RegFilePlugin_regFile[12][22] , \RegFilePlugin_regFile[12][21] ,
         \RegFilePlugin_regFile[12][20] , \RegFilePlugin_regFile[12][19] ,
         \RegFilePlugin_regFile[12][18] , \RegFilePlugin_regFile[12][17] ,
         \RegFilePlugin_regFile[12][16] , \RegFilePlugin_regFile[12][15] ,
         \RegFilePlugin_regFile[12][14] , \RegFilePlugin_regFile[12][13] ,
         \RegFilePlugin_regFile[12][12] , \RegFilePlugin_regFile[12][11] ,
         \RegFilePlugin_regFile[12][10] , \RegFilePlugin_regFile[12][9] ,
         \RegFilePlugin_regFile[12][8] , \RegFilePlugin_regFile[12][7] ,
         \RegFilePlugin_regFile[12][6] , \RegFilePlugin_regFile[12][5] ,
         \RegFilePlugin_regFile[12][4] , \RegFilePlugin_regFile[12][3] ,
         \RegFilePlugin_regFile[12][2] , \RegFilePlugin_regFile[12][1] ,
         \RegFilePlugin_regFile[12][0] , \RegFilePlugin_regFile[13][31] ,
         \RegFilePlugin_regFile[13][30] , \RegFilePlugin_regFile[13][29] ,
         \RegFilePlugin_regFile[13][28] , \RegFilePlugin_regFile[13][27] ,
         \RegFilePlugin_regFile[13][26] , \RegFilePlugin_regFile[13][25] ,
         \RegFilePlugin_regFile[13][24] , \RegFilePlugin_regFile[13][23] ,
         \RegFilePlugin_regFile[13][22] , \RegFilePlugin_regFile[13][21] ,
         \RegFilePlugin_regFile[13][20] , \RegFilePlugin_regFile[13][19] ,
         \RegFilePlugin_regFile[13][18] , \RegFilePlugin_regFile[13][17] ,
         \RegFilePlugin_regFile[13][16] , \RegFilePlugin_regFile[13][15] ,
         \RegFilePlugin_regFile[13][14] , \RegFilePlugin_regFile[13][13] ,
         \RegFilePlugin_regFile[13][12] , \RegFilePlugin_regFile[13][11] ,
         \RegFilePlugin_regFile[13][10] , \RegFilePlugin_regFile[13][9] ,
         \RegFilePlugin_regFile[13][8] , \RegFilePlugin_regFile[13][7] ,
         \RegFilePlugin_regFile[13][6] , \RegFilePlugin_regFile[13][5] ,
         \RegFilePlugin_regFile[13][4] , \RegFilePlugin_regFile[13][3] ,
         \RegFilePlugin_regFile[13][2] , \RegFilePlugin_regFile[13][1] ,
         \RegFilePlugin_regFile[13][0] , \RegFilePlugin_regFile[14][31] ,
         \RegFilePlugin_regFile[14][30] , \RegFilePlugin_regFile[14][29] ,
         \RegFilePlugin_regFile[14][28] , \RegFilePlugin_regFile[14][27] ,
         \RegFilePlugin_regFile[14][26] , \RegFilePlugin_regFile[14][25] ,
         \RegFilePlugin_regFile[14][24] , \RegFilePlugin_regFile[14][23] ,
         \RegFilePlugin_regFile[14][22] , \RegFilePlugin_regFile[14][21] ,
         \RegFilePlugin_regFile[14][20] , \RegFilePlugin_regFile[14][19] ,
         \RegFilePlugin_regFile[14][18] , \RegFilePlugin_regFile[14][17] ,
         \RegFilePlugin_regFile[14][16] , \RegFilePlugin_regFile[14][15] ,
         \RegFilePlugin_regFile[14][14] , \RegFilePlugin_regFile[14][13] ,
         \RegFilePlugin_regFile[14][12] , \RegFilePlugin_regFile[14][11] ,
         \RegFilePlugin_regFile[14][10] , \RegFilePlugin_regFile[14][9] ,
         \RegFilePlugin_regFile[14][8] , \RegFilePlugin_regFile[14][7] ,
         \RegFilePlugin_regFile[14][6] , \RegFilePlugin_regFile[14][5] ,
         \RegFilePlugin_regFile[14][4] , \RegFilePlugin_regFile[14][3] ,
         \RegFilePlugin_regFile[14][2] , \RegFilePlugin_regFile[14][1] ,
         \RegFilePlugin_regFile[14][0] , \RegFilePlugin_regFile[15][31] ,
         \RegFilePlugin_regFile[15][30] , \RegFilePlugin_regFile[15][29] ,
         \RegFilePlugin_regFile[15][28] , \RegFilePlugin_regFile[15][27] ,
         \RegFilePlugin_regFile[15][26] , \RegFilePlugin_regFile[15][25] ,
         \RegFilePlugin_regFile[15][24] , \RegFilePlugin_regFile[15][23] ,
         \RegFilePlugin_regFile[15][22] , \RegFilePlugin_regFile[15][21] ,
         \RegFilePlugin_regFile[15][20] , \RegFilePlugin_regFile[15][19] ,
         \RegFilePlugin_regFile[15][18] , \RegFilePlugin_regFile[15][17] ,
         \RegFilePlugin_regFile[15][16] , \RegFilePlugin_regFile[15][15] ,
         \RegFilePlugin_regFile[15][14] , \RegFilePlugin_regFile[15][13] ,
         \RegFilePlugin_regFile[15][12] , \RegFilePlugin_regFile[15][11] ,
         \RegFilePlugin_regFile[15][10] , \RegFilePlugin_regFile[15][9] ,
         \RegFilePlugin_regFile[15][8] , \RegFilePlugin_regFile[15][7] ,
         \RegFilePlugin_regFile[15][6] , \RegFilePlugin_regFile[15][5] ,
         \RegFilePlugin_regFile[15][4] , \RegFilePlugin_regFile[15][3] ,
         \RegFilePlugin_regFile[15][2] , \RegFilePlugin_regFile[15][1] ,
         \RegFilePlugin_regFile[15][0] , \RegFilePlugin_regFile[16][31] ,
         \RegFilePlugin_regFile[16][30] , \RegFilePlugin_regFile[16][29] ,
         \RegFilePlugin_regFile[16][28] , \RegFilePlugin_regFile[16][27] ,
         \RegFilePlugin_regFile[16][26] , \RegFilePlugin_regFile[16][25] ,
         \RegFilePlugin_regFile[16][24] , \RegFilePlugin_regFile[16][23] ,
         \RegFilePlugin_regFile[16][22] , \RegFilePlugin_regFile[16][21] ,
         \RegFilePlugin_regFile[16][20] , \RegFilePlugin_regFile[16][19] ,
         \RegFilePlugin_regFile[16][18] , \RegFilePlugin_regFile[16][17] ,
         \RegFilePlugin_regFile[16][16] , \RegFilePlugin_regFile[16][15] ,
         \RegFilePlugin_regFile[16][14] , \RegFilePlugin_regFile[16][13] ,
         \RegFilePlugin_regFile[16][12] , \RegFilePlugin_regFile[16][11] ,
         \RegFilePlugin_regFile[16][10] , \RegFilePlugin_regFile[16][9] ,
         \RegFilePlugin_regFile[16][8] , \RegFilePlugin_regFile[16][7] ,
         \RegFilePlugin_regFile[16][6] , \RegFilePlugin_regFile[16][5] ,
         \RegFilePlugin_regFile[16][4] , \RegFilePlugin_regFile[16][3] ,
         \RegFilePlugin_regFile[16][2] , \RegFilePlugin_regFile[16][1] ,
         \RegFilePlugin_regFile[16][0] , \RegFilePlugin_regFile[17][31] ,
         \RegFilePlugin_regFile[17][30] , \RegFilePlugin_regFile[17][29] ,
         \RegFilePlugin_regFile[17][28] , \RegFilePlugin_regFile[17][27] ,
         \RegFilePlugin_regFile[17][26] , \RegFilePlugin_regFile[17][25] ,
         \RegFilePlugin_regFile[17][24] , \RegFilePlugin_regFile[17][23] ,
         \RegFilePlugin_regFile[17][22] , \RegFilePlugin_regFile[17][21] ,
         \RegFilePlugin_regFile[17][20] , \RegFilePlugin_regFile[17][19] ,
         \RegFilePlugin_regFile[17][18] , \RegFilePlugin_regFile[17][17] ,
         \RegFilePlugin_regFile[17][16] , \RegFilePlugin_regFile[17][15] ,
         \RegFilePlugin_regFile[17][14] , \RegFilePlugin_regFile[17][13] ,
         \RegFilePlugin_regFile[17][12] , \RegFilePlugin_regFile[17][11] ,
         \RegFilePlugin_regFile[17][10] , \RegFilePlugin_regFile[17][9] ,
         \RegFilePlugin_regFile[17][8] , \RegFilePlugin_regFile[17][7] ,
         \RegFilePlugin_regFile[17][6] , \RegFilePlugin_regFile[17][5] ,
         \RegFilePlugin_regFile[17][4] , \RegFilePlugin_regFile[17][3] ,
         \RegFilePlugin_regFile[17][2] , \RegFilePlugin_regFile[17][1] ,
         \RegFilePlugin_regFile[17][0] , \RegFilePlugin_regFile[18][31] ,
         \RegFilePlugin_regFile[18][30] , \RegFilePlugin_regFile[18][29] ,
         \RegFilePlugin_regFile[18][28] , \RegFilePlugin_regFile[18][27] ,
         \RegFilePlugin_regFile[18][26] , \RegFilePlugin_regFile[18][25] ,
         \RegFilePlugin_regFile[18][24] , \RegFilePlugin_regFile[18][23] ,
         \RegFilePlugin_regFile[18][22] , \RegFilePlugin_regFile[18][21] ,
         \RegFilePlugin_regFile[18][20] , \RegFilePlugin_regFile[18][19] ,
         \RegFilePlugin_regFile[18][18] , \RegFilePlugin_regFile[18][17] ,
         \RegFilePlugin_regFile[18][16] , \RegFilePlugin_regFile[18][15] ,
         \RegFilePlugin_regFile[18][14] , \RegFilePlugin_regFile[18][13] ,
         \RegFilePlugin_regFile[18][12] , \RegFilePlugin_regFile[18][11] ,
         \RegFilePlugin_regFile[18][10] , \RegFilePlugin_regFile[18][9] ,
         \RegFilePlugin_regFile[18][8] , \RegFilePlugin_regFile[18][7] ,
         \RegFilePlugin_regFile[18][6] , \RegFilePlugin_regFile[18][5] ,
         \RegFilePlugin_regFile[18][4] , \RegFilePlugin_regFile[18][3] ,
         \RegFilePlugin_regFile[18][2] , \RegFilePlugin_regFile[18][1] ,
         \RegFilePlugin_regFile[18][0] , \RegFilePlugin_regFile[19][31] ,
         \RegFilePlugin_regFile[19][30] , \RegFilePlugin_regFile[19][29] ,
         \RegFilePlugin_regFile[19][28] , \RegFilePlugin_regFile[19][27] ,
         \RegFilePlugin_regFile[19][26] , \RegFilePlugin_regFile[19][25] ,
         \RegFilePlugin_regFile[19][24] , \RegFilePlugin_regFile[19][23] ,
         \RegFilePlugin_regFile[19][22] , \RegFilePlugin_regFile[19][21] ,
         \RegFilePlugin_regFile[19][20] , \RegFilePlugin_regFile[19][19] ,
         \RegFilePlugin_regFile[19][18] , \RegFilePlugin_regFile[19][17] ,
         \RegFilePlugin_regFile[19][16] , \RegFilePlugin_regFile[19][15] ,
         \RegFilePlugin_regFile[19][14] , \RegFilePlugin_regFile[19][13] ,
         \RegFilePlugin_regFile[19][12] , \RegFilePlugin_regFile[19][11] ,
         \RegFilePlugin_regFile[19][10] , \RegFilePlugin_regFile[19][9] ,
         \RegFilePlugin_regFile[19][8] , \RegFilePlugin_regFile[19][7] ,
         \RegFilePlugin_regFile[19][6] , \RegFilePlugin_regFile[19][5] ,
         \RegFilePlugin_regFile[19][4] , \RegFilePlugin_regFile[19][3] ,
         \RegFilePlugin_regFile[19][2] , \RegFilePlugin_regFile[19][1] ,
         \RegFilePlugin_regFile[19][0] , \RegFilePlugin_regFile[20][31] ,
         \RegFilePlugin_regFile[20][30] , \RegFilePlugin_regFile[20][29] ,
         \RegFilePlugin_regFile[20][28] , \RegFilePlugin_regFile[20][27] ,
         \RegFilePlugin_regFile[20][26] , \RegFilePlugin_regFile[20][25] ,
         \RegFilePlugin_regFile[20][24] , \RegFilePlugin_regFile[20][23] ,
         \RegFilePlugin_regFile[20][22] , \RegFilePlugin_regFile[20][21] ,
         \RegFilePlugin_regFile[20][20] , \RegFilePlugin_regFile[20][19] ,
         \RegFilePlugin_regFile[20][18] , \RegFilePlugin_regFile[20][17] ,
         \RegFilePlugin_regFile[20][16] , \RegFilePlugin_regFile[20][15] ,
         \RegFilePlugin_regFile[20][14] , \RegFilePlugin_regFile[20][13] ,
         \RegFilePlugin_regFile[20][12] , \RegFilePlugin_regFile[20][11] ,
         \RegFilePlugin_regFile[20][10] , \RegFilePlugin_regFile[20][9] ,
         \RegFilePlugin_regFile[20][8] , \RegFilePlugin_regFile[20][7] ,
         \RegFilePlugin_regFile[20][6] , \RegFilePlugin_regFile[20][5] ,
         \RegFilePlugin_regFile[20][4] , \RegFilePlugin_regFile[20][3] ,
         \RegFilePlugin_regFile[20][2] , \RegFilePlugin_regFile[20][1] ,
         \RegFilePlugin_regFile[20][0] , \RegFilePlugin_regFile[21][31] ,
         \RegFilePlugin_regFile[21][30] , \RegFilePlugin_regFile[21][29] ,
         \RegFilePlugin_regFile[21][28] , \RegFilePlugin_regFile[21][27] ,
         \RegFilePlugin_regFile[21][26] , \RegFilePlugin_regFile[21][25] ,
         \RegFilePlugin_regFile[21][24] , \RegFilePlugin_regFile[21][23] ,
         \RegFilePlugin_regFile[21][22] , \RegFilePlugin_regFile[21][21] ,
         \RegFilePlugin_regFile[21][20] , \RegFilePlugin_regFile[21][19] ,
         \RegFilePlugin_regFile[21][18] , \RegFilePlugin_regFile[21][17] ,
         \RegFilePlugin_regFile[21][16] , \RegFilePlugin_regFile[21][15] ,
         \RegFilePlugin_regFile[21][14] , \RegFilePlugin_regFile[21][13] ,
         \RegFilePlugin_regFile[21][12] , \RegFilePlugin_regFile[21][11] ,
         \RegFilePlugin_regFile[21][10] , \RegFilePlugin_regFile[21][9] ,
         \RegFilePlugin_regFile[21][8] , \RegFilePlugin_regFile[21][7] ,
         \RegFilePlugin_regFile[21][6] , \RegFilePlugin_regFile[21][5] ,
         \RegFilePlugin_regFile[21][4] , \RegFilePlugin_regFile[21][3] ,
         \RegFilePlugin_regFile[21][2] , \RegFilePlugin_regFile[21][1] ,
         \RegFilePlugin_regFile[21][0] , \RegFilePlugin_regFile[22][31] ,
         \RegFilePlugin_regFile[22][30] , \RegFilePlugin_regFile[22][29] ,
         \RegFilePlugin_regFile[22][28] , \RegFilePlugin_regFile[22][27] ,
         \RegFilePlugin_regFile[22][26] , \RegFilePlugin_regFile[22][25] ,
         \RegFilePlugin_regFile[22][24] , \RegFilePlugin_regFile[22][23] ,
         \RegFilePlugin_regFile[22][22] , \RegFilePlugin_regFile[22][21] ,
         \RegFilePlugin_regFile[22][20] , \RegFilePlugin_regFile[22][19] ,
         \RegFilePlugin_regFile[22][18] , \RegFilePlugin_regFile[22][17] ,
         \RegFilePlugin_regFile[22][16] , \RegFilePlugin_regFile[22][15] ,
         \RegFilePlugin_regFile[22][14] , \RegFilePlugin_regFile[22][13] ,
         \RegFilePlugin_regFile[22][12] , \RegFilePlugin_regFile[22][11] ,
         \RegFilePlugin_regFile[22][10] , \RegFilePlugin_regFile[22][9] ,
         \RegFilePlugin_regFile[22][8] , \RegFilePlugin_regFile[22][7] ,
         \RegFilePlugin_regFile[22][6] , \RegFilePlugin_regFile[22][5] ,
         \RegFilePlugin_regFile[22][4] , \RegFilePlugin_regFile[22][3] ,
         \RegFilePlugin_regFile[22][2] , \RegFilePlugin_regFile[22][1] ,
         \RegFilePlugin_regFile[22][0] , \RegFilePlugin_regFile[23][31] ,
         \RegFilePlugin_regFile[23][30] , \RegFilePlugin_regFile[23][29] ,
         \RegFilePlugin_regFile[23][28] , \RegFilePlugin_regFile[23][27] ,
         \RegFilePlugin_regFile[23][26] , \RegFilePlugin_regFile[23][25] ,
         \RegFilePlugin_regFile[23][24] , \RegFilePlugin_regFile[23][23] ,
         \RegFilePlugin_regFile[23][22] , \RegFilePlugin_regFile[23][21] ,
         \RegFilePlugin_regFile[23][20] , \RegFilePlugin_regFile[23][19] ,
         \RegFilePlugin_regFile[23][18] , \RegFilePlugin_regFile[23][17] ,
         \RegFilePlugin_regFile[23][16] , \RegFilePlugin_regFile[23][15] ,
         \RegFilePlugin_regFile[23][14] , \RegFilePlugin_regFile[23][13] ,
         \RegFilePlugin_regFile[23][12] , \RegFilePlugin_regFile[23][11] ,
         \RegFilePlugin_regFile[23][10] , \RegFilePlugin_regFile[23][9] ,
         \RegFilePlugin_regFile[23][8] , \RegFilePlugin_regFile[23][7] ,
         \RegFilePlugin_regFile[23][6] , \RegFilePlugin_regFile[23][5] ,
         \RegFilePlugin_regFile[23][4] , \RegFilePlugin_regFile[23][3] ,
         \RegFilePlugin_regFile[23][2] , \RegFilePlugin_regFile[23][1] ,
         \RegFilePlugin_regFile[23][0] , \RegFilePlugin_regFile[24][31] ,
         \RegFilePlugin_regFile[24][30] , \RegFilePlugin_regFile[24][29] ,
         \RegFilePlugin_regFile[24][28] , \RegFilePlugin_regFile[24][27] ,
         \RegFilePlugin_regFile[24][26] , \RegFilePlugin_regFile[24][25] ,
         \RegFilePlugin_regFile[24][24] , \RegFilePlugin_regFile[24][23] ,
         \RegFilePlugin_regFile[24][22] , \RegFilePlugin_regFile[24][21] ,
         \RegFilePlugin_regFile[24][20] , \RegFilePlugin_regFile[24][19] ,
         \RegFilePlugin_regFile[24][18] , \RegFilePlugin_regFile[24][17] ,
         \RegFilePlugin_regFile[24][16] , \RegFilePlugin_regFile[24][15] ,
         \RegFilePlugin_regFile[24][14] , \RegFilePlugin_regFile[24][13] ,
         \RegFilePlugin_regFile[24][12] , \RegFilePlugin_regFile[24][11] ,
         \RegFilePlugin_regFile[24][10] , \RegFilePlugin_regFile[24][9] ,
         \RegFilePlugin_regFile[24][8] , \RegFilePlugin_regFile[24][7] ,
         \RegFilePlugin_regFile[24][6] , \RegFilePlugin_regFile[24][5] ,
         \RegFilePlugin_regFile[24][4] , \RegFilePlugin_regFile[24][3] ,
         \RegFilePlugin_regFile[24][2] , \RegFilePlugin_regFile[24][1] ,
         \RegFilePlugin_regFile[24][0] , \RegFilePlugin_regFile[25][31] ,
         \RegFilePlugin_regFile[25][30] , \RegFilePlugin_regFile[25][29] ,
         \RegFilePlugin_regFile[25][28] , \RegFilePlugin_regFile[25][27] ,
         \RegFilePlugin_regFile[25][26] , \RegFilePlugin_regFile[25][25] ,
         \RegFilePlugin_regFile[25][24] , \RegFilePlugin_regFile[25][23] ,
         \RegFilePlugin_regFile[25][22] , \RegFilePlugin_regFile[25][21] ,
         \RegFilePlugin_regFile[25][20] , \RegFilePlugin_regFile[25][19] ,
         \RegFilePlugin_regFile[25][18] , \RegFilePlugin_regFile[25][17] ,
         \RegFilePlugin_regFile[25][16] , \RegFilePlugin_regFile[25][15] ,
         \RegFilePlugin_regFile[25][14] , \RegFilePlugin_regFile[25][13] ,
         \RegFilePlugin_regFile[25][12] , \RegFilePlugin_regFile[25][11] ,
         \RegFilePlugin_regFile[25][10] , \RegFilePlugin_regFile[25][9] ,
         \RegFilePlugin_regFile[25][8] , \RegFilePlugin_regFile[25][7] ,
         \RegFilePlugin_regFile[25][6] , \RegFilePlugin_regFile[25][5] ,
         \RegFilePlugin_regFile[25][4] , \RegFilePlugin_regFile[25][3] ,
         \RegFilePlugin_regFile[25][2] , \RegFilePlugin_regFile[25][1] ,
         \RegFilePlugin_regFile[25][0] , \RegFilePlugin_regFile[26][31] ,
         \RegFilePlugin_regFile[26][30] , \RegFilePlugin_regFile[26][29] ,
         \RegFilePlugin_regFile[26][28] , \RegFilePlugin_regFile[26][27] ,
         \RegFilePlugin_regFile[26][26] , \RegFilePlugin_regFile[26][25] ,
         \RegFilePlugin_regFile[26][24] , \RegFilePlugin_regFile[26][23] ,
         \RegFilePlugin_regFile[26][22] , \RegFilePlugin_regFile[26][21] ,
         \RegFilePlugin_regFile[26][20] , \RegFilePlugin_regFile[26][19] ,
         \RegFilePlugin_regFile[26][18] , \RegFilePlugin_regFile[26][17] ,
         \RegFilePlugin_regFile[26][16] , \RegFilePlugin_regFile[26][15] ,
         \RegFilePlugin_regFile[26][14] , \RegFilePlugin_regFile[26][13] ,
         \RegFilePlugin_regFile[26][12] , \RegFilePlugin_regFile[26][11] ,
         \RegFilePlugin_regFile[26][10] , \RegFilePlugin_regFile[26][9] ,
         \RegFilePlugin_regFile[26][8] , \RegFilePlugin_regFile[26][7] ,
         \RegFilePlugin_regFile[26][6] , \RegFilePlugin_regFile[26][5] ,
         \RegFilePlugin_regFile[26][4] , \RegFilePlugin_regFile[26][3] ,
         \RegFilePlugin_regFile[26][2] , \RegFilePlugin_regFile[26][1] ,
         \RegFilePlugin_regFile[26][0] , \RegFilePlugin_regFile[27][31] ,
         \RegFilePlugin_regFile[27][30] , \RegFilePlugin_regFile[27][29] ,
         \RegFilePlugin_regFile[27][28] , \RegFilePlugin_regFile[27][27] ,
         \RegFilePlugin_regFile[27][26] , \RegFilePlugin_regFile[27][25] ,
         \RegFilePlugin_regFile[27][24] , \RegFilePlugin_regFile[27][23] ,
         \RegFilePlugin_regFile[27][22] , \RegFilePlugin_regFile[27][21] ,
         \RegFilePlugin_regFile[27][20] , \RegFilePlugin_regFile[27][19] ,
         \RegFilePlugin_regFile[27][18] , \RegFilePlugin_regFile[27][17] ,
         \RegFilePlugin_regFile[27][16] , \RegFilePlugin_regFile[27][15] ,
         \RegFilePlugin_regFile[27][14] , \RegFilePlugin_regFile[27][13] ,
         \RegFilePlugin_regFile[27][12] , \RegFilePlugin_regFile[27][11] ,
         \RegFilePlugin_regFile[27][10] , \RegFilePlugin_regFile[27][9] ,
         \RegFilePlugin_regFile[27][8] , \RegFilePlugin_regFile[27][7] ,
         \RegFilePlugin_regFile[27][6] , \RegFilePlugin_regFile[27][5] ,
         \RegFilePlugin_regFile[27][4] , \RegFilePlugin_regFile[27][3] ,
         \RegFilePlugin_regFile[27][2] , \RegFilePlugin_regFile[27][1] ,
         \RegFilePlugin_regFile[27][0] , \RegFilePlugin_regFile[28][31] ,
         \RegFilePlugin_regFile[28][30] , \RegFilePlugin_regFile[28][29] ,
         \RegFilePlugin_regFile[28][28] , \RegFilePlugin_regFile[28][27] ,
         \RegFilePlugin_regFile[28][26] , \RegFilePlugin_regFile[28][25] ,
         \RegFilePlugin_regFile[28][24] , \RegFilePlugin_regFile[28][23] ,
         \RegFilePlugin_regFile[28][22] , \RegFilePlugin_regFile[28][21] ,
         \RegFilePlugin_regFile[28][20] , \RegFilePlugin_regFile[28][19] ,
         \RegFilePlugin_regFile[28][18] , \RegFilePlugin_regFile[28][17] ,
         \RegFilePlugin_regFile[28][16] , \RegFilePlugin_regFile[28][15] ,
         \RegFilePlugin_regFile[28][14] , \RegFilePlugin_regFile[28][13] ,
         \RegFilePlugin_regFile[28][12] , \RegFilePlugin_regFile[28][11] ,
         \RegFilePlugin_regFile[28][10] , \RegFilePlugin_regFile[28][9] ,
         \RegFilePlugin_regFile[28][8] , \RegFilePlugin_regFile[28][7] ,
         \RegFilePlugin_regFile[28][6] , \RegFilePlugin_regFile[28][5] ,
         \RegFilePlugin_regFile[28][4] , \RegFilePlugin_regFile[28][3] ,
         \RegFilePlugin_regFile[28][2] , \RegFilePlugin_regFile[28][1] ,
         \RegFilePlugin_regFile[28][0] , \RegFilePlugin_regFile[29][31] ,
         \RegFilePlugin_regFile[29][30] , \RegFilePlugin_regFile[29][29] ,
         \RegFilePlugin_regFile[29][28] , \RegFilePlugin_regFile[29][27] ,
         \RegFilePlugin_regFile[29][26] , \RegFilePlugin_regFile[29][25] ,
         \RegFilePlugin_regFile[29][24] , \RegFilePlugin_regFile[29][23] ,
         \RegFilePlugin_regFile[29][22] , \RegFilePlugin_regFile[29][21] ,
         \RegFilePlugin_regFile[29][20] , \RegFilePlugin_regFile[29][19] ,
         \RegFilePlugin_regFile[29][18] , \RegFilePlugin_regFile[29][17] ,
         \RegFilePlugin_regFile[29][16] , \RegFilePlugin_regFile[29][15] ,
         \RegFilePlugin_regFile[29][14] , \RegFilePlugin_regFile[29][13] ,
         \RegFilePlugin_regFile[29][12] , \RegFilePlugin_regFile[29][11] ,
         \RegFilePlugin_regFile[29][10] , \RegFilePlugin_regFile[29][9] ,
         \RegFilePlugin_regFile[29][8] , \RegFilePlugin_regFile[29][7] ,
         \RegFilePlugin_regFile[29][6] , \RegFilePlugin_regFile[29][5] ,
         \RegFilePlugin_regFile[29][4] , \RegFilePlugin_regFile[29][3] ,
         \RegFilePlugin_regFile[29][2] , \RegFilePlugin_regFile[29][1] ,
         \RegFilePlugin_regFile[29][0] , \RegFilePlugin_regFile[30][31] ,
         \RegFilePlugin_regFile[30][30] , \RegFilePlugin_regFile[30][29] ,
         \RegFilePlugin_regFile[30][28] , \RegFilePlugin_regFile[30][27] ,
         \RegFilePlugin_regFile[30][26] , \RegFilePlugin_regFile[30][25] ,
         \RegFilePlugin_regFile[30][24] , \RegFilePlugin_regFile[30][23] ,
         \RegFilePlugin_regFile[30][22] , \RegFilePlugin_regFile[30][21] ,
         \RegFilePlugin_regFile[30][20] , \RegFilePlugin_regFile[30][19] ,
         \RegFilePlugin_regFile[30][18] , \RegFilePlugin_regFile[30][17] ,
         \RegFilePlugin_regFile[30][16] , \RegFilePlugin_regFile[30][15] ,
         \RegFilePlugin_regFile[30][14] , \RegFilePlugin_regFile[30][13] ,
         \RegFilePlugin_regFile[30][12] , \RegFilePlugin_regFile[30][11] ,
         \RegFilePlugin_regFile[30][10] , \RegFilePlugin_regFile[30][9] ,
         \RegFilePlugin_regFile[30][8] , \RegFilePlugin_regFile[30][7] ,
         \RegFilePlugin_regFile[30][6] , \RegFilePlugin_regFile[30][5] ,
         \RegFilePlugin_regFile[30][4] , \RegFilePlugin_regFile[30][3] ,
         \RegFilePlugin_regFile[30][2] , \RegFilePlugin_regFile[30][1] ,
         \RegFilePlugin_regFile[30][0] , \RegFilePlugin_regFile[31][31] ,
         \RegFilePlugin_regFile[31][30] , \RegFilePlugin_regFile[31][29] ,
         \RegFilePlugin_regFile[31][28] , \RegFilePlugin_regFile[31][27] ,
         \RegFilePlugin_regFile[31][26] , \RegFilePlugin_regFile[31][25] ,
         \RegFilePlugin_regFile[31][24] , \RegFilePlugin_regFile[31][23] ,
         \RegFilePlugin_regFile[31][22] , \RegFilePlugin_regFile[31][21] ,
         \RegFilePlugin_regFile[31][20] , \RegFilePlugin_regFile[31][19] ,
         \RegFilePlugin_regFile[31][18] , \RegFilePlugin_regFile[31][17] ,
         \RegFilePlugin_regFile[31][16] , \RegFilePlugin_regFile[31][15] ,
         \RegFilePlugin_regFile[31][14] , \RegFilePlugin_regFile[31][13] ,
         \RegFilePlugin_regFile[31][12] , \RegFilePlugin_regFile[31][11] ,
         \RegFilePlugin_regFile[31][10] , \RegFilePlugin_regFile[31][9] ,
         \RegFilePlugin_regFile[31][8] , \RegFilePlugin_regFile[31][7] ,
         \RegFilePlugin_regFile[31][6] , \RegFilePlugin_regFile[31][5] ,
         \RegFilePlugin_regFile[31][4] , \RegFilePlugin_regFile[31][3] ,
         \RegFilePlugin_regFile[31][2] , \RegFilePlugin_regFile[31][1] ,
         \RegFilePlugin_regFile[31][0] , N823, N824, N825, N826, N827, N828,
         N829, N830, N831, N832, N833, N834, N835, N836, N837, N838, N839,
         N840, N841, N842, N843, N844, N845, N846, N847, N848, N849, N850,
         N851, N852, N853, N854, N856, N857, N858, N859, N860, N861, N862,
         N863, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873,
         N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884,
         N885, N886, N887, iBus_rsp_valid, DebugPlugin_haltIt,
         execute_DO_EBREAK, execute_CSR_WRITE_OPCODE, execute_IS_CSR,
         memory_BRANCH_DO, execute_REGFILE_WRITE_VALID,
         memory_REGFILE_WRITE_VALID, memory_INSTRUCTION_29,
         memory_INSTRUCTION_28, writeBack_REGFILE_WRITE_VALID,
         execute_SRC_LESS_UNSIGNED, execute_SRC2_FORCE_ZERO,
         _zz_lastStageRegFileWrite_payload_address_29,
         _zz_lastStageRegFileWrite_payload_address_28, writeBack_MEMORY_ENABLE,
         memory_ALIGNEMENT_FAULT, memory_MEMORY_ENABLE, execute_MEMORY_ENABLE,
         lastStageIsValid, DebugPlugin_godmode,
         IBusCachedPlugin_fetchPc_booted,
         _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1,
         IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid,
         execute_arbitration_isValid, memory_arbitration_isValid,
         execute_LightShifterPlugin_isActive,
         HazardSimplePlugin_writeBackBuffer_valid, CsrPlugin_mie_MTIE,
         CsrPlugin_mip_MSIP, CsrPlugin_mie_MSIE, CsrPlugin_mip_MEIP,
         CsrPlugin_mie_MEIE, CsrPlugin_exceptionPendings_0,
         CsrPlugin_exceptionPendings_1, CsrPlugin_exceptionPendings_2,
         CsrPlugin_exceptionPendings_3, CsrPlugin_mstatus_MIE,
         CsrPlugin_interrupt_valid, CsrPlugin_hadException,
         CsrPlugin_pipelineLiberator_pcValids_2, \CsrPlugin_interrupt_code[3] ,
         execute_CsrPlugin_csr_768, execute_CsrPlugin_csr_836,
         execute_CsrPlugin_csr_772, execute_CsrPlugin_csr_773,
         execute_CsrPlugin_csr_833, execute_CsrPlugin_csr_834,
         execute_CsrPlugin_csr_835, execute_CsrPlugin_csr_3008,
         execute_CsrPlugin_csr_4032, DebugPlugin_isPipBusy,
         DebugPlugin_debugUsed, DebugPlugin_disableEbreak, DebugPlugin_resetIt,
         DebugPlugin_haltedByBreak, DebugPlugin_stepIt,
         _zz_when_DebugPlugin_l244, CsrPlugin_mstatus_MPIE,
         CsrPlugin_mcause_interrupt, when_InstructionCache_l239,
         CsrPlugin_pipelineLiberator_pcValids_0,
         CsrPlugin_pipelineLiberator_pcValids_1, N1771, N1781, N1782, N1783,
         N1784, N1785, N1792, N1840, N2007, N2076, N2210,
         \IBusCachedPlugin_cache/decodeStage_hit_valid ,
         \IBusCachedPlugin_cache/lineLoader_cmdSent ,
         \IBusCachedPlugin_cache/_zz_when_InstructionCache_l342 ,
         \IBusCachedPlugin_cache/lineLoader_flushCounter[0] ,
         \IBusCachedPlugin_cache/lineLoader_flushPending ,
         \IBusCachedPlugin_cache/lineLoader_valid ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[27] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[26] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[25] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[24] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[23] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[22] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[21] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[20] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[19] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[18] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[17] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[16] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[15] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[14] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[13] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[12] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[11] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[10] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[9] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[8] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[7] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[6] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[5] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[4] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[3] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[2] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[0] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][27] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][26] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][25] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][24] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][23] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][22] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][21] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][20] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][19] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][18] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][17] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][16] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][15] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][14] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][13] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][12] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][11] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][10] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][9] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][8] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][7] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][6] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][5] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][4] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][3] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][2] ,
         \IBusCachedPlugin_cache/ways_0_tags[0][0] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][27] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][26] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][25] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][24] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][23] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][22] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][21] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][20] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][19] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][18] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][17] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][16] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][15] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][14] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][13] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][12] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][11] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][10] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][9] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][8] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][7] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][6] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][5] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][4] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][3] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][2] ,
         \IBusCachedPlugin_cache/ways_0_tags[1][0] ,
         \IBusCachedPlugin_cache/banks_0[0][31] ,
         \IBusCachedPlugin_cache/banks_0[0][30] ,
         \IBusCachedPlugin_cache/banks_0[0][29] ,
         \IBusCachedPlugin_cache/banks_0[0][28] ,
         \IBusCachedPlugin_cache/banks_0[0][27] ,
         \IBusCachedPlugin_cache/banks_0[0][26] ,
         \IBusCachedPlugin_cache/banks_0[0][25] ,
         \IBusCachedPlugin_cache/banks_0[0][24] ,
         \IBusCachedPlugin_cache/banks_0[0][23] ,
         \IBusCachedPlugin_cache/banks_0[0][22] ,
         \IBusCachedPlugin_cache/banks_0[0][21] ,
         \IBusCachedPlugin_cache/banks_0[0][20] ,
         \IBusCachedPlugin_cache/banks_0[0][19] ,
         \IBusCachedPlugin_cache/banks_0[0][18] ,
         \IBusCachedPlugin_cache/banks_0[0][17] ,
         \IBusCachedPlugin_cache/banks_0[0][16] ,
         \IBusCachedPlugin_cache/banks_0[0][15] ,
         \IBusCachedPlugin_cache/banks_0[0][14] ,
         \IBusCachedPlugin_cache/banks_0[0][13] ,
         \IBusCachedPlugin_cache/banks_0[0][12] ,
         \IBusCachedPlugin_cache/banks_0[0][11] ,
         \IBusCachedPlugin_cache/banks_0[0][10] ,
         \IBusCachedPlugin_cache/banks_0[0][9] ,
         \IBusCachedPlugin_cache/banks_0[0][8] ,
         \IBusCachedPlugin_cache/banks_0[0][7] ,
         \IBusCachedPlugin_cache/banks_0[0][6] ,
         \IBusCachedPlugin_cache/banks_0[0][5] ,
         \IBusCachedPlugin_cache/banks_0[0][4] ,
         \IBusCachedPlugin_cache/banks_0[0][3] ,
         \IBusCachedPlugin_cache/banks_0[0][2] ,
         \IBusCachedPlugin_cache/banks_0[0][1] ,
         \IBusCachedPlugin_cache/banks_0[0][0] ,
         \IBusCachedPlugin_cache/banks_0[1][31] ,
         \IBusCachedPlugin_cache/banks_0[1][30] ,
         \IBusCachedPlugin_cache/banks_0[1][29] ,
         \IBusCachedPlugin_cache/banks_0[1][28] ,
         \IBusCachedPlugin_cache/banks_0[1][27] ,
         \IBusCachedPlugin_cache/banks_0[1][26] ,
         \IBusCachedPlugin_cache/banks_0[1][25] ,
         \IBusCachedPlugin_cache/banks_0[1][24] ,
         \IBusCachedPlugin_cache/banks_0[1][23] ,
         \IBusCachedPlugin_cache/banks_0[1][22] ,
         \IBusCachedPlugin_cache/banks_0[1][21] ,
         \IBusCachedPlugin_cache/banks_0[1][20] ,
         \IBusCachedPlugin_cache/banks_0[1][19] ,
         \IBusCachedPlugin_cache/banks_0[1][18] ,
         \IBusCachedPlugin_cache/banks_0[1][17] ,
         \IBusCachedPlugin_cache/banks_0[1][16] ,
         \IBusCachedPlugin_cache/banks_0[1][15] ,
         \IBusCachedPlugin_cache/banks_0[1][14] ,
         \IBusCachedPlugin_cache/banks_0[1][13] ,
         \IBusCachedPlugin_cache/banks_0[1][12] ,
         \IBusCachedPlugin_cache/banks_0[1][11] ,
         \IBusCachedPlugin_cache/banks_0[1][10] ,
         \IBusCachedPlugin_cache/banks_0[1][9] ,
         \IBusCachedPlugin_cache/banks_0[1][8] ,
         \IBusCachedPlugin_cache/banks_0[1][7] ,
         \IBusCachedPlugin_cache/banks_0[1][6] ,
         \IBusCachedPlugin_cache/banks_0[1][5] ,
         \IBusCachedPlugin_cache/banks_0[1][4] ,
         \IBusCachedPlugin_cache/banks_0[1][3] ,
         \IBusCachedPlugin_cache/banks_0[1][2] ,
         \IBusCachedPlugin_cache/banks_0[1][1] ,
         \IBusCachedPlugin_cache/banks_0[1][0] ,
         \IBusCachedPlugin_cache/banks_0[2][31] ,
         \IBusCachedPlugin_cache/banks_0[2][30] ,
         \IBusCachedPlugin_cache/banks_0[2][29] ,
         \IBusCachedPlugin_cache/banks_0[2][28] ,
         \IBusCachedPlugin_cache/banks_0[2][27] ,
         \IBusCachedPlugin_cache/banks_0[2][26] ,
         \IBusCachedPlugin_cache/banks_0[2][25] ,
         \IBusCachedPlugin_cache/banks_0[2][24] ,
         \IBusCachedPlugin_cache/banks_0[2][23] ,
         \IBusCachedPlugin_cache/banks_0[2][22] ,
         \IBusCachedPlugin_cache/banks_0[2][21] ,
         \IBusCachedPlugin_cache/banks_0[2][20] ,
         \IBusCachedPlugin_cache/banks_0[2][19] ,
         \IBusCachedPlugin_cache/banks_0[2][18] ,
         \IBusCachedPlugin_cache/banks_0[2][17] ,
         \IBusCachedPlugin_cache/banks_0[2][16] ,
         \IBusCachedPlugin_cache/banks_0[2][15] ,
         \IBusCachedPlugin_cache/banks_0[2][14] ,
         \IBusCachedPlugin_cache/banks_0[2][13] ,
         \IBusCachedPlugin_cache/banks_0[2][12] ,
         \IBusCachedPlugin_cache/banks_0[2][11] ,
         \IBusCachedPlugin_cache/banks_0[2][10] ,
         \IBusCachedPlugin_cache/banks_0[2][9] ,
         \IBusCachedPlugin_cache/banks_0[2][8] ,
         \IBusCachedPlugin_cache/banks_0[2][7] ,
         \IBusCachedPlugin_cache/banks_0[2][6] ,
         \IBusCachedPlugin_cache/banks_0[2][5] ,
         \IBusCachedPlugin_cache/banks_0[2][4] ,
         \IBusCachedPlugin_cache/banks_0[2][3] ,
         \IBusCachedPlugin_cache/banks_0[2][2] ,
         \IBusCachedPlugin_cache/banks_0[2][1] ,
         \IBusCachedPlugin_cache/banks_0[2][0] ,
         \IBusCachedPlugin_cache/banks_0[3][31] ,
         \IBusCachedPlugin_cache/banks_0[3][30] ,
         \IBusCachedPlugin_cache/banks_0[3][29] ,
         \IBusCachedPlugin_cache/banks_0[3][28] ,
         \IBusCachedPlugin_cache/banks_0[3][27] ,
         \IBusCachedPlugin_cache/banks_0[3][26] ,
         \IBusCachedPlugin_cache/banks_0[3][25] ,
         \IBusCachedPlugin_cache/banks_0[3][24] ,
         \IBusCachedPlugin_cache/banks_0[3][23] ,
         \IBusCachedPlugin_cache/banks_0[3][22] ,
         \IBusCachedPlugin_cache/banks_0[3][21] ,
         \IBusCachedPlugin_cache/banks_0[3][20] ,
         \IBusCachedPlugin_cache/banks_0[3][19] ,
         \IBusCachedPlugin_cache/banks_0[3][18] ,
         \IBusCachedPlugin_cache/banks_0[3][17] ,
         \IBusCachedPlugin_cache/banks_0[3][16] ,
         \IBusCachedPlugin_cache/banks_0[3][15] ,
         \IBusCachedPlugin_cache/banks_0[3][14] ,
         \IBusCachedPlugin_cache/banks_0[3][13] ,
         \IBusCachedPlugin_cache/banks_0[3][12] ,
         \IBusCachedPlugin_cache/banks_0[3][11] ,
         \IBusCachedPlugin_cache/banks_0[3][10] ,
         \IBusCachedPlugin_cache/banks_0[3][9] ,
         \IBusCachedPlugin_cache/banks_0[3][8] ,
         \IBusCachedPlugin_cache/banks_0[3][7] ,
         \IBusCachedPlugin_cache/banks_0[3][6] ,
         \IBusCachedPlugin_cache/banks_0[3][5] ,
         \IBusCachedPlugin_cache/banks_0[3][4] ,
         \IBusCachedPlugin_cache/banks_0[3][3] ,
         \IBusCachedPlugin_cache/banks_0[3][2] ,
         \IBusCachedPlugin_cache/banks_0[3][1] ,
         \IBusCachedPlugin_cache/banks_0[3][0] ,
         \IBusCachedPlugin_cache/banks_0[4][31] ,
         \IBusCachedPlugin_cache/banks_0[4][30] ,
         \IBusCachedPlugin_cache/banks_0[4][29] ,
         \IBusCachedPlugin_cache/banks_0[4][28] ,
         \IBusCachedPlugin_cache/banks_0[4][27] ,
         \IBusCachedPlugin_cache/banks_0[4][26] ,
         \IBusCachedPlugin_cache/banks_0[4][25] ,
         \IBusCachedPlugin_cache/banks_0[4][24] ,
         \IBusCachedPlugin_cache/banks_0[4][23] ,
         \IBusCachedPlugin_cache/banks_0[4][22] ,
         \IBusCachedPlugin_cache/banks_0[4][21] ,
         \IBusCachedPlugin_cache/banks_0[4][20] ,
         \IBusCachedPlugin_cache/banks_0[4][19] ,
         \IBusCachedPlugin_cache/banks_0[4][18] ,
         \IBusCachedPlugin_cache/banks_0[4][17] ,
         \IBusCachedPlugin_cache/banks_0[4][16] ,
         \IBusCachedPlugin_cache/banks_0[4][15] ,
         \IBusCachedPlugin_cache/banks_0[4][14] ,
         \IBusCachedPlugin_cache/banks_0[4][13] ,
         \IBusCachedPlugin_cache/banks_0[4][12] ,
         \IBusCachedPlugin_cache/banks_0[4][11] ,
         \IBusCachedPlugin_cache/banks_0[4][10] ,
         \IBusCachedPlugin_cache/banks_0[4][9] ,
         \IBusCachedPlugin_cache/banks_0[4][8] ,
         \IBusCachedPlugin_cache/banks_0[4][7] ,
         \IBusCachedPlugin_cache/banks_0[4][6] ,
         \IBusCachedPlugin_cache/banks_0[4][5] ,
         \IBusCachedPlugin_cache/banks_0[4][4] ,
         \IBusCachedPlugin_cache/banks_0[4][3] ,
         \IBusCachedPlugin_cache/banks_0[4][2] ,
         \IBusCachedPlugin_cache/banks_0[4][1] ,
         \IBusCachedPlugin_cache/banks_0[4][0] ,
         \IBusCachedPlugin_cache/banks_0[5][31] ,
         \IBusCachedPlugin_cache/banks_0[5][30] ,
         \IBusCachedPlugin_cache/banks_0[5][29] ,
         \IBusCachedPlugin_cache/banks_0[5][28] ,
         \IBusCachedPlugin_cache/banks_0[5][27] ,
         \IBusCachedPlugin_cache/banks_0[5][26] ,
         \IBusCachedPlugin_cache/banks_0[5][25] ,
         \IBusCachedPlugin_cache/banks_0[5][24] ,
         \IBusCachedPlugin_cache/banks_0[5][23] ,
         \IBusCachedPlugin_cache/banks_0[5][22] ,
         \IBusCachedPlugin_cache/banks_0[5][21] ,
         \IBusCachedPlugin_cache/banks_0[5][20] ,
         \IBusCachedPlugin_cache/banks_0[5][19] ,
         \IBusCachedPlugin_cache/banks_0[5][18] ,
         \IBusCachedPlugin_cache/banks_0[5][17] ,
         \IBusCachedPlugin_cache/banks_0[5][16] ,
         \IBusCachedPlugin_cache/banks_0[5][15] ,
         \IBusCachedPlugin_cache/banks_0[5][14] ,
         \IBusCachedPlugin_cache/banks_0[5][13] ,
         \IBusCachedPlugin_cache/banks_0[5][12] ,
         \IBusCachedPlugin_cache/banks_0[5][11] ,
         \IBusCachedPlugin_cache/banks_0[5][10] ,
         \IBusCachedPlugin_cache/banks_0[5][9] ,
         \IBusCachedPlugin_cache/banks_0[5][8] ,
         \IBusCachedPlugin_cache/banks_0[5][7] ,
         \IBusCachedPlugin_cache/banks_0[5][6] ,
         \IBusCachedPlugin_cache/banks_0[5][5] ,
         \IBusCachedPlugin_cache/banks_0[5][4] ,
         \IBusCachedPlugin_cache/banks_0[5][3] ,
         \IBusCachedPlugin_cache/banks_0[5][2] ,
         \IBusCachedPlugin_cache/banks_0[5][1] ,
         \IBusCachedPlugin_cache/banks_0[5][0] ,
         \IBusCachedPlugin_cache/banks_0[6][31] ,
         \IBusCachedPlugin_cache/banks_0[6][30] ,
         \IBusCachedPlugin_cache/banks_0[6][29] ,
         \IBusCachedPlugin_cache/banks_0[6][28] ,
         \IBusCachedPlugin_cache/banks_0[6][27] ,
         \IBusCachedPlugin_cache/banks_0[6][26] ,
         \IBusCachedPlugin_cache/banks_0[6][25] ,
         \IBusCachedPlugin_cache/banks_0[6][24] ,
         \IBusCachedPlugin_cache/banks_0[6][23] ,
         \IBusCachedPlugin_cache/banks_0[6][22] ,
         \IBusCachedPlugin_cache/banks_0[6][21] ,
         \IBusCachedPlugin_cache/banks_0[6][20] ,
         \IBusCachedPlugin_cache/banks_0[6][19] ,
         \IBusCachedPlugin_cache/banks_0[6][18] ,
         \IBusCachedPlugin_cache/banks_0[6][17] ,
         \IBusCachedPlugin_cache/banks_0[6][16] ,
         \IBusCachedPlugin_cache/banks_0[6][15] ,
         \IBusCachedPlugin_cache/banks_0[6][14] ,
         \IBusCachedPlugin_cache/banks_0[6][13] ,
         \IBusCachedPlugin_cache/banks_0[6][12] ,
         \IBusCachedPlugin_cache/banks_0[6][11] ,
         \IBusCachedPlugin_cache/banks_0[6][10] ,
         \IBusCachedPlugin_cache/banks_0[6][9] ,
         \IBusCachedPlugin_cache/banks_0[6][8] ,
         \IBusCachedPlugin_cache/banks_0[6][7] ,
         \IBusCachedPlugin_cache/banks_0[6][6] ,
         \IBusCachedPlugin_cache/banks_0[6][5] ,
         \IBusCachedPlugin_cache/banks_0[6][4] ,
         \IBusCachedPlugin_cache/banks_0[6][3] ,
         \IBusCachedPlugin_cache/banks_0[6][2] ,
         \IBusCachedPlugin_cache/banks_0[6][1] ,
         \IBusCachedPlugin_cache/banks_0[6][0] ,
         \IBusCachedPlugin_cache/banks_0[7][31] ,
         \IBusCachedPlugin_cache/banks_0[7][30] ,
         \IBusCachedPlugin_cache/banks_0[7][29] ,
         \IBusCachedPlugin_cache/banks_0[7][28] ,
         \IBusCachedPlugin_cache/banks_0[7][27] ,
         \IBusCachedPlugin_cache/banks_0[7][26] ,
         \IBusCachedPlugin_cache/banks_0[7][25] ,
         \IBusCachedPlugin_cache/banks_0[7][24] ,
         \IBusCachedPlugin_cache/banks_0[7][23] ,
         \IBusCachedPlugin_cache/banks_0[7][22] ,
         \IBusCachedPlugin_cache/banks_0[7][21] ,
         \IBusCachedPlugin_cache/banks_0[7][20] ,
         \IBusCachedPlugin_cache/banks_0[7][19] ,
         \IBusCachedPlugin_cache/banks_0[7][18] ,
         \IBusCachedPlugin_cache/banks_0[7][17] ,
         \IBusCachedPlugin_cache/banks_0[7][16] ,
         \IBusCachedPlugin_cache/banks_0[7][15] ,
         \IBusCachedPlugin_cache/banks_0[7][14] ,
         \IBusCachedPlugin_cache/banks_0[7][13] ,
         \IBusCachedPlugin_cache/banks_0[7][12] ,
         \IBusCachedPlugin_cache/banks_0[7][11] ,
         \IBusCachedPlugin_cache/banks_0[7][10] ,
         \IBusCachedPlugin_cache/banks_0[7][9] ,
         \IBusCachedPlugin_cache/banks_0[7][8] ,
         \IBusCachedPlugin_cache/banks_0[7][7] ,
         \IBusCachedPlugin_cache/banks_0[7][6] ,
         \IBusCachedPlugin_cache/banks_0[7][5] ,
         \IBusCachedPlugin_cache/banks_0[7][4] ,
         \IBusCachedPlugin_cache/banks_0[7][3] ,
         \IBusCachedPlugin_cache/banks_0[7][2] ,
         \IBusCachedPlugin_cache/banks_0[7][1] ,
         \IBusCachedPlugin_cache/banks_0[7][0] ,
         \IBusCachedPlugin_cache/banks_0[8][31] ,
         \IBusCachedPlugin_cache/banks_0[8][30] ,
         \IBusCachedPlugin_cache/banks_0[8][29] ,
         \IBusCachedPlugin_cache/banks_0[8][28] ,
         \IBusCachedPlugin_cache/banks_0[8][27] ,
         \IBusCachedPlugin_cache/banks_0[8][26] ,
         \IBusCachedPlugin_cache/banks_0[8][25] ,
         \IBusCachedPlugin_cache/banks_0[8][24] ,
         \IBusCachedPlugin_cache/banks_0[8][23] ,
         \IBusCachedPlugin_cache/banks_0[8][22] ,
         \IBusCachedPlugin_cache/banks_0[8][21] ,
         \IBusCachedPlugin_cache/banks_0[8][20] ,
         \IBusCachedPlugin_cache/banks_0[8][19] ,
         \IBusCachedPlugin_cache/banks_0[8][18] ,
         \IBusCachedPlugin_cache/banks_0[8][17] ,
         \IBusCachedPlugin_cache/banks_0[8][16] ,
         \IBusCachedPlugin_cache/banks_0[8][15] ,
         \IBusCachedPlugin_cache/banks_0[8][14] ,
         \IBusCachedPlugin_cache/banks_0[8][13] ,
         \IBusCachedPlugin_cache/banks_0[8][12] ,
         \IBusCachedPlugin_cache/banks_0[8][11] ,
         \IBusCachedPlugin_cache/banks_0[8][10] ,
         \IBusCachedPlugin_cache/banks_0[8][9] ,
         \IBusCachedPlugin_cache/banks_0[8][8] ,
         \IBusCachedPlugin_cache/banks_0[8][7] ,
         \IBusCachedPlugin_cache/banks_0[8][6] ,
         \IBusCachedPlugin_cache/banks_0[8][5] ,
         \IBusCachedPlugin_cache/banks_0[8][4] ,
         \IBusCachedPlugin_cache/banks_0[8][3] ,
         \IBusCachedPlugin_cache/banks_0[8][2] ,
         \IBusCachedPlugin_cache/banks_0[8][1] ,
         \IBusCachedPlugin_cache/banks_0[8][0] ,
         \IBusCachedPlugin_cache/banks_0[9][31] ,
         \IBusCachedPlugin_cache/banks_0[9][30] ,
         \IBusCachedPlugin_cache/banks_0[9][29] ,
         \IBusCachedPlugin_cache/banks_0[9][28] ,
         \IBusCachedPlugin_cache/banks_0[9][27] ,
         \IBusCachedPlugin_cache/banks_0[9][26] ,
         \IBusCachedPlugin_cache/banks_0[9][25] ,
         \IBusCachedPlugin_cache/banks_0[9][24] ,
         \IBusCachedPlugin_cache/banks_0[9][23] ,
         \IBusCachedPlugin_cache/banks_0[9][22] ,
         \IBusCachedPlugin_cache/banks_0[9][21] ,
         \IBusCachedPlugin_cache/banks_0[9][20] ,
         \IBusCachedPlugin_cache/banks_0[9][19] ,
         \IBusCachedPlugin_cache/banks_0[9][18] ,
         \IBusCachedPlugin_cache/banks_0[9][17] ,
         \IBusCachedPlugin_cache/banks_0[9][16] ,
         \IBusCachedPlugin_cache/banks_0[9][15] ,
         \IBusCachedPlugin_cache/banks_0[9][14] ,
         \IBusCachedPlugin_cache/banks_0[9][13] ,
         \IBusCachedPlugin_cache/banks_0[9][12] ,
         \IBusCachedPlugin_cache/banks_0[9][11] ,
         \IBusCachedPlugin_cache/banks_0[9][10] ,
         \IBusCachedPlugin_cache/banks_0[9][9] ,
         \IBusCachedPlugin_cache/banks_0[9][8] ,
         \IBusCachedPlugin_cache/banks_0[9][7] ,
         \IBusCachedPlugin_cache/banks_0[9][6] ,
         \IBusCachedPlugin_cache/banks_0[9][5] ,
         \IBusCachedPlugin_cache/banks_0[9][4] ,
         \IBusCachedPlugin_cache/banks_0[9][3] ,
         \IBusCachedPlugin_cache/banks_0[9][2] ,
         \IBusCachedPlugin_cache/banks_0[9][1] ,
         \IBusCachedPlugin_cache/banks_0[9][0] ,
         \IBusCachedPlugin_cache/banks_0[10][31] ,
         \IBusCachedPlugin_cache/banks_0[10][30] ,
         \IBusCachedPlugin_cache/banks_0[10][29] ,
         \IBusCachedPlugin_cache/banks_0[10][28] ,
         \IBusCachedPlugin_cache/banks_0[10][27] ,
         \IBusCachedPlugin_cache/banks_0[10][26] ,
         \IBusCachedPlugin_cache/banks_0[10][25] ,
         \IBusCachedPlugin_cache/banks_0[10][24] ,
         \IBusCachedPlugin_cache/banks_0[10][23] ,
         \IBusCachedPlugin_cache/banks_0[10][22] ,
         \IBusCachedPlugin_cache/banks_0[10][21] ,
         \IBusCachedPlugin_cache/banks_0[10][20] ,
         \IBusCachedPlugin_cache/banks_0[10][19] ,
         \IBusCachedPlugin_cache/banks_0[10][18] ,
         \IBusCachedPlugin_cache/banks_0[10][17] ,
         \IBusCachedPlugin_cache/banks_0[10][16] ,
         \IBusCachedPlugin_cache/banks_0[10][15] ,
         \IBusCachedPlugin_cache/banks_0[10][14] ,
         \IBusCachedPlugin_cache/banks_0[10][13] ,
         \IBusCachedPlugin_cache/banks_0[10][12] ,
         \IBusCachedPlugin_cache/banks_0[10][11] ,
         \IBusCachedPlugin_cache/banks_0[10][10] ,
         \IBusCachedPlugin_cache/banks_0[10][9] ,
         \IBusCachedPlugin_cache/banks_0[10][8] ,
         \IBusCachedPlugin_cache/banks_0[10][7] ,
         \IBusCachedPlugin_cache/banks_0[10][6] ,
         \IBusCachedPlugin_cache/banks_0[10][5] ,
         \IBusCachedPlugin_cache/banks_0[10][4] ,
         \IBusCachedPlugin_cache/banks_0[10][3] ,
         \IBusCachedPlugin_cache/banks_0[10][2] ,
         \IBusCachedPlugin_cache/banks_0[10][1] ,
         \IBusCachedPlugin_cache/banks_0[10][0] ,
         \IBusCachedPlugin_cache/banks_0[11][31] ,
         \IBusCachedPlugin_cache/banks_0[11][30] ,
         \IBusCachedPlugin_cache/banks_0[11][29] ,
         \IBusCachedPlugin_cache/banks_0[11][28] ,
         \IBusCachedPlugin_cache/banks_0[11][27] ,
         \IBusCachedPlugin_cache/banks_0[11][26] ,
         \IBusCachedPlugin_cache/banks_0[11][25] ,
         \IBusCachedPlugin_cache/banks_0[11][24] ,
         \IBusCachedPlugin_cache/banks_0[11][23] ,
         \IBusCachedPlugin_cache/banks_0[11][22] ,
         \IBusCachedPlugin_cache/banks_0[11][21] ,
         \IBusCachedPlugin_cache/banks_0[11][20] ,
         \IBusCachedPlugin_cache/banks_0[11][19] ,
         \IBusCachedPlugin_cache/banks_0[11][18] ,
         \IBusCachedPlugin_cache/banks_0[11][17] ,
         \IBusCachedPlugin_cache/banks_0[11][16] ,
         \IBusCachedPlugin_cache/banks_0[11][15] ,
         \IBusCachedPlugin_cache/banks_0[11][14] ,
         \IBusCachedPlugin_cache/banks_0[11][13] ,
         \IBusCachedPlugin_cache/banks_0[11][12] ,
         \IBusCachedPlugin_cache/banks_0[11][11] ,
         \IBusCachedPlugin_cache/banks_0[11][10] ,
         \IBusCachedPlugin_cache/banks_0[11][9] ,
         \IBusCachedPlugin_cache/banks_0[11][8] ,
         \IBusCachedPlugin_cache/banks_0[11][7] ,
         \IBusCachedPlugin_cache/banks_0[11][6] ,
         \IBusCachedPlugin_cache/banks_0[11][5] ,
         \IBusCachedPlugin_cache/banks_0[11][4] ,
         \IBusCachedPlugin_cache/banks_0[11][3] ,
         \IBusCachedPlugin_cache/banks_0[11][2] ,
         \IBusCachedPlugin_cache/banks_0[11][1] ,
         \IBusCachedPlugin_cache/banks_0[11][0] ,
         \IBusCachedPlugin_cache/banks_0[12][31] ,
         \IBusCachedPlugin_cache/banks_0[12][30] ,
         \IBusCachedPlugin_cache/banks_0[12][29] ,
         \IBusCachedPlugin_cache/banks_0[12][28] ,
         \IBusCachedPlugin_cache/banks_0[12][27] ,
         \IBusCachedPlugin_cache/banks_0[12][26] ,
         \IBusCachedPlugin_cache/banks_0[12][25] ,
         \IBusCachedPlugin_cache/banks_0[12][24] ,
         \IBusCachedPlugin_cache/banks_0[12][23] ,
         \IBusCachedPlugin_cache/banks_0[12][22] ,
         \IBusCachedPlugin_cache/banks_0[12][21] ,
         \IBusCachedPlugin_cache/banks_0[12][20] ,
         \IBusCachedPlugin_cache/banks_0[12][19] ,
         \IBusCachedPlugin_cache/banks_0[12][18] ,
         \IBusCachedPlugin_cache/banks_0[12][17] ,
         \IBusCachedPlugin_cache/banks_0[12][16] ,
         \IBusCachedPlugin_cache/banks_0[12][15] ,
         \IBusCachedPlugin_cache/banks_0[12][14] ,
         \IBusCachedPlugin_cache/banks_0[12][13] ,
         \IBusCachedPlugin_cache/banks_0[12][12] ,
         \IBusCachedPlugin_cache/banks_0[12][11] ,
         \IBusCachedPlugin_cache/banks_0[12][10] ,
         \IBusCachedPlugin_cache/banks_0[12][9] ,
         \IBusCachedPlugin_cache/banks_0[12][8] ,
         \IBusCachedPlugin_cache/banks_0[12][7] ,
         \IBusCachedPlugin_cache/banks_0[12][6] ,
         \IBusCachedPlugin_cache/banks_0[12][5] ,
         \IBusCachedPlugin_cache/banks_0[12][4] ,
         \IBusCachedPlugin_cache/banks_0[12][3] ,
         \IBusCachedPlugin_cache/banks_0[12][2] ,
         \IBusCachedPlugin_cache/banks_0[12][1] ,
         \IBusCachedPlugin_cache/banks_0[12][0] ,
         \IBusCachedPlugin_cache/banks_0[13][31] ,
         \IBusCachedPlugin_cache/banks_0[13][30] ,
         \IBusCachedPlugin_cache/banks_0[13][29] ,
         \IBusCachedPlugin_cache/banks_0[13][28] ,
         \IBusCachedPlugin_cache/banks_0[13][27] ,
         \IBusCachedPlugin_cache/banks_0[13][26] ,
         \IBusCachedPlugin_cache/banks_0[13][25] ,
         \IBusCachedPlugin_cache/banks_0[13][24] ,
         \IBusCachedPlugin_cache/banks_0[13][23] ,
         \IBusCachedPlugin_cache/banks_0[13][22] ,
         \IBusCachedPlugin_cache/banks_0[13][21] ,
         \IBusCachedPlugin_cache/banks_0[13][20] ,
         \IBusCachedPlugin_cache/banks_0[13][19] ,
         \IBusCachedPlugin_cache/banks_0[13][18] ,
         \IBusCachedPlugin_cache/banks_0[13][17] ,
         \IBusCachedPlugin_cache/banks_0[13][16] ,
         \IBusCachedPlugin_cache/banks_0[13][15] ,
         \IBusCachedPlugin_cache/banks_0[13][14] ,
         \IBusCachedPlugin_cache/banks_0[13][13] ,
         \IBusCachedPlugin_cache/banks_0[13][12] ,
         \IBusCachedPlugin_cache/banks_0[13][11] ,
         \IBusCachedPlugin_cache/banks_0[13][10] ,
         \IBusCachedPlugin_cache/banks_0[13][9] ,
         \IBusCachedPlugin_cache/banks_0[13][8] ,
         \IBusCachedPlugin_cache/banks_0[13][7] ,
         \IBusCachedPlugin_cache/banks_0[13][6] ,
         \IBusCachedPlugin_cache/banks_0[13][5] ,
         \IBusCachedPlugin_cache/banks_0[13][4] ,
         \IBusCachedPlugin_cache/banks_0[13][3] ,
         \IBusCachedPlugin_cache/banks_0[13][2] ,
         \IBusCachedPlugin_cache/banks_0[13][1] ,
         \IBusCachedPlugin_cache/banks_0[13][0] ,
         \IBusCachedPlugin_cache/banks_0[14][31] ,
         \IBusCachedPlugin_cache/banks_0[14][30] ,
         \IBusCachedPlugin_cache/banks_0[14][29] ,
         \IBusCachedPlugin_cache/banks_0[14][28] ,
         \IBusCachedPlugin_cache/banks_0[14][27] ,
         \IBusCachedPlugin_cache/banks_0[14][26] ,
         \IBusCachedPlugin_cache/banks_0[14][25] ,
         \IBusCachedPlugin_cache/banks_0[14][24] ,
         \IBusCachedPlugin_cache/banks_0[14][23] ,
         \IBusCachedPlugin_cache/banks_0[14][22] ,
         \IBusCachedPlugin_cache/banks_0[14][21] ,
         \IBusCachedPlugin_cache/banks_0[14][20] ,
         \IBusCachedPlugin_cache/banks_0[14][19] ,
         \IBusCachedPlugin_cache/banks_0[14][18] ,
         \IBusCachedPlugin_cache/banks_0[14][17] ,
         \IBusCachedPlugin_cache/banks_0[14][16] ,
         \IBusCachedPlugin_cache/banks_0[14][15] ,
         \IBusCachedPlugin_cache/banks_0[14][14] ,
         \IBusCachedPlugin_cache/banks_0[14][13] ,
         \IBusCachedPlugin_cache/banks_0[14][12] ,
         \IBusCachedPlugin_cache/banks_0[14][11] ,
         \IBusCachedPlugin_cache/banks_0[14][10] ,
         \IBusCachedPlugin_cache/banks_0[14][9] ,
         \IBusCachedPlugin_cache/banks_0[14][8] ,
         \IBusCachedPlugin_cache/banks_0[14][7] ,
         \IBusCachedPlugin_cache/banks_0[14][6] ,
         \IBusCachedPlugin_cache/banks_0[14][5] ,
         \IBusCachedPlugin_cache/banks_0[14][4] ,
         \IBusCachedPlugin_cache/banks_0[14][3] ,
         \IBusCachedPlugin_cache/banks_0[14][2] ,
         \IBusCachedPlugin_cache/banks_0[14][1] ,
         \IBusCachedPlugin_cache/banks_0[14][0] ,
         \IBusCachedPlugin_cache/banks_0[15][31] ,
         \IBusCachedPlugin_cache/banks_0[15][30] ,
         \IBusCachedPlugin_cache/banks_0[15][29] ,
         \IBusCachedPlugin_cache/banks_0[15][28] ,
         \IBusCachedPlugin_cache/banks_0[15][27] ,
         \IBusCachedPlugin_cache/banks_0[15][26] ,
         \IBusCachedPlugin_cache/banks_0[15][25] ,
         \IBusCachedPlugin_cache/banks_0[15][24] ,
         \IBusCachedPlugin_cache/banks_0[15][23] ,
         \IBusCachedPlugin_cache/banks_0[15][22] ,
         \IBusCachedPlugin_cache/banks_0[15][21] ,
         \IBusCachedPlugin_cache/banks_0[15][20] ,
         \IBusCachedPlugin_cache/banks_0[15][19] ,
         \IBusCachedPlugin_cache/banks_0[15][18] ,
         \IBusCachedPlugin_cache/banks_0[15][17] ,
         \IBusCachedPlugin_cache/banks_0[15][16] ,
         \IBusCachedPlugin_cache/banks_0[15][15] ,
         \IBusCachedPlugin_cache/banks_0[15][14] ,
         \IBusCachedPlugin_cache/banks_0[15][13] ,
         \IBusCachedPlugin_cache/banks_0[15][12] ,
         \IBusCachedPlugin_cache/banks_0[15][11] ,
         \IBusCachedPlugin_cache/banks_0[15][10] ,
         \IBusCachedPlugin_cache/banks_0[15][9] ,
         \IBusCachedPlugin_cache/banks_0[15][8] ,
         \IBusCachedPlugin_cache/banks_0[15][7] ,
         \IBusCachedPlugin_cache/banks_0[15][6] ,
         \IBusCachedPlugin_cache/banks_0[15][5] ,
         \IBusCachedPlugin_cache/banks_0[15][4] ,
         \IBusCachedPlugin_cache/banks_0[15][3] ,
         \IBusCachedPlugin_cache/banks_0[15][2] ,
         \IBusCachedPlugin_cache/banks_0[15][1] ,
         \IBusCachedPlugin_cache/banks_0[15][0] ,
         \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[2] ,
         \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[1] ,
         \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[0] ,
         \IBusCachedPlugin_cache/_zz_ways_0_tags_port[0] ,
         \IBusCachedPlugin_cache/n23 , \IBusCachedPlugin_cache/n22 ,
         \IBusCachedPlugin_cache/n21 , \IBusCachedPlugin_cache/n20 ,
         \IBusCachedPlugin_cache/n19 , \IBusCachedPlugin_cache/n18 ,
         \IBusCachedPlugin_cache/n17 , \IBusCachedPlugin_cache/n16 ,
         \IBusCachedPlugin_cache/n15 , \IBusCachedPlugin_cache/n14 ,
         \IBusCachedPlugin_cache/n13 , \IBusCachedPlugin_cache/n12 ,
         \IBusCachedPlugin_cache/n11 , \IBusCachedPlugin_cache/n10 ,
         \IBusCachedPlugin_cache/n9 , \IBusCachedPlugin_cache/n8 ,
         \IBusCachedPlugin_cache/n7 , \IBusCachedPlugin_cache/n6 ,
         \IBusCachedPlugin_cache/n5 , \IBusCachedPlugin_cache/n4 ,
         \IBusCachedPlugin_cache/n3 , \IBusCachedPlugin_cache/n2 , n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4023, n4024, n4025, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n4022, n4026, n4061, n4079, n5319, n5320, n5321, n5322,
         n5323, n6121, n6122, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264;
  wire   [29:0] iBusWishbone_ADR;
  wire   [4:0] _zz__zz_execute_SRC1_1;
  wire   [6:0] execute_INSTRUCTION;
  wire   [11:0] _zz__zz_execute_SRC2_3;
  wire   [1:0] execute_SHIFT_CTRL;
  wire   [13:10] _zz__zz_execute_BranchPlugin_branch_src2;
  wire   [19:15] decode_INSTRUCTION;
  wire   [6:0] _zz_decode_LEGAL_INSTRUCTION_1;
  wire   [29:25] _zz_decode_LEGAL_INSTRUCTION_13;
  wire   [31:0] _zz_RegFilePlugin_regFile_port0;
  wire   [31:0] _zz_RegFilePlugin_regFile_port1;
  wire   [31:0] IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  wire   [31:0] IBusCachedPlugin_cache_io_cpu_fetch_data;
  wire   [31:0] IBusCachedPlugin_cache_io_cpu_decode_physicalAddress;
  wire   [31:0] iBus_rsp_payload_data;
  wire   [2:0] switch_Fetcher_l362;
  wire   [31:0] writeBack_REGFILE_WRITE_DATA;
  wire   [1:0] memory_MEMORY_ADDRESS_LOW;
  wire   [31:0] memory_PC;
  wire   [1:0] memory_ENV_CTRL;
  wire   [1:0] execute_ENV_CTRL;
  wire   [1:0] writeBack_ENV_CTRL;
  wire   [31:0] memory_BRANCH_CALC;
  wire   [31:0] execute_PC;
  wire   [31:0] execute_RS1;
  wire   [1:0] execute_BRANCH_CTRL;
  wire   [14:7] memory_INSTRUCTION;
  wire   [1:0] execute_SRC2_CTRL;
  wire   [1:0] execute_SRC1_CTRL;
  wire   [1:0] execute_ALU_CTRL;
  wire   [1:0] execute_ALU_BITWISE_CTRL;
  wire   [14:7] _zz_lastStageRegFileWrite_payload_address;
  wire   [1:0] writeBack_MEMORY_ADDRESS_LOW;
  wire   [31:0] memory_REGFILE_WRITE_DATA;
  wire   [31:0] execute_RS2;
  wire   [31:0] writeBack_PC;
  wire   [31:0] CsrPlugin_mepc;
  wire   [31:0] IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  wire   [4:0] execute_LightShifterPlugin_amplitudeReg;
  wire   [4:0] HazardSimplePlugin_writeBackBuffer_payload_address;
  wire   [3:0] CsrPlugin_exceptionPortCtrl_exceptionContext_code;
  wire   [29:0] CsrPlugin_mtvec_base;
  wire   [31:0] _zz_CsrPlugin_csrMapping_readDataInit;
  wire   [31:0] externalInterruptArray_regNext;
  wire   [4:0] DebugPlugin_busReadDataReg;
  wire   [1:0] CsrPlugin_mstatus_MPP;
  wire   [3:0] CsrPlugin_mcause_exceptionCode;
  wire   [31:0] CsrPlugin_mtval;
  wire   [1:0] dBus_cmd_halfPipe_payload_address;
  wire   [1:0] dBus_cmd_halfPipe_payload_size;
  wire   [31:0] CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr;
  assign \iBusWishbone_ADR[29]  = iBusWishbone_ADR[29];
  assign \iBusWishbone_ADR[28]  = iBusWishbone_ADR[28];
  assign \iBusWishbone_ADR[27]  = iBusWishbone_ADR[27];
  assign \iBusWishbone_ADR[26]  = iBusWishbone_ADR[26];
  assign \iBusWishbone_ADR[25]  = iBusWishbone_ADR[25];
  assign \iBusWishbone_ADR[24]  = iBusWishbone_ADR[24];
  assign \iBusWishbone_ADR[23]  = iBusWishbone_ADR[23];
  assign \iBusWishbone_ADR[22]  = iBusWishbone_ADR[22];
  assign \iBusWishbone_ADR[21]  = iBusWishbone_ADR[21];
  assign \iBusWishbone_ADR[20]  = iBusWishbone_ADR[20];
  assign \iBusWishbone_ADR[19]  = iBusWishbone_ADR[19];
  assign \iBusWishbone_ADR[18]  = iBusWishbone_ADR[18];
  assign \iBusWishbone_ADR[17]  = iBusWishbone_ADR[17];
  assign \iBusWishbone_ADR[16]  = iBusWishbone_ADR[16];
  assign \iBusWishbone_ADR[15]  = iBusWishbone_ADR[15];
  assign \iBusWishbone_ADR[14]  = iBusWishbone_ADR[14];
  assign \iBusWishbone_ADR[13]  = iBusWishbone_ADR[13];
  assign \iBusWishbone_ADR[12]  = iBusWishbone_ADR[12];
  assign \iBusWishbone_ADR[11]  = iBusWishbone_ADR[11];
  assign \iBusWishbone_ADR[10]  = iBusWishbone_ADR[10];
  assign \iBusWishbone_ADR[9]  = iBusWishbone_ADR[9];
  assign \iBusWishbone_ADR[8]  = iBusWishbone_ADR[8];
  assign \iBusWishbone_ADR[7]  = iBusWishbone_ADR[7];
  assign \iBusWishbone_ADR[6]  = iBusWishbone_ADR[6];
  assign \iBusWishbone_ADR[5]  = iBusWishbone_ADR[5];
  assign \iBusWishbone_ADR[4]  = iBusWishbone_ADR[4];
  assign \iBusWishbone_ADR[2]  = iBusWishbone_ADR[2];
  assign \iBusWishbone_ADR[1]  = iBusWishbone_ADR[1];
  assign \iBusWishbone_ADR[0]  = iBusWishbone_ADR[0];
  assign iBusWishbone_CYC = when_InstructionCache_l239;

  dfnrq1 IBusCachedPlugin_fetchPc_booted_reg ( .D(n7121), .CP(n7252), .Q(
        IBusCachedPlugin_fetchPc_booted) );
  dfnrq1 \externalInterruptArray_regNext_reg[7]  ( .D(
        externalInterruptArray[7]), .CP(n7252), .Q(
        externalInterruptArray_regNext[7]) );
  dfnrq1 \externalInterruptArray_regNext_reg[6]  ( .D(
        externalInterruptArray[6]), .CP(n7224), .Q(
        externalInterruptArray_regNext[6]) );
  dfnrq1 \externalInterruptArray_regNext_reg[5]  ( .D(
        externalInterruptArray[5]), .CP(n7252), .Q(
        externalInterruptArray_regNext[5]) );
  dfnrq1 \externalInterruptArray_regNext_reg[4]  ( .D(
        externalInterruptArray[4]), .CP(n7231), .Q(
        externalInterruptArray_regNext[4]) );
  dfnrq1 \externalInterruptArray_regNext_reg[3]  ( .D(
        externalInterruptArray[3]), .CP(n7224), .Q(
        externalInterruptArray_regNext[3]) );
  dfnrq1 \externalInterruptArray_regNext_reg[2]  ( .D(
        externalInterruptArray[2]), .CP(n7224), .Q(
        externalInterruptArray_regNext[2]) );
  dfnrq1 \externalInterruptArray_regNext_reg[1]  ( .D(
        externalInterruptArray[1]), .CP(n7222), .Q(
        externalInterruptArray_regNext[1]) );
  dfnrq1 \externalInterruptArray_regNext_reg[0]  ( .D(
        externalInterruptArray[0]), .CP(n7223), .Q(
        externalInterruptArray_regNext[0]) );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[31]  ( .D(
        iBusWishbone_DAT_MISO[31]), .CP(n7225), .Q(iBus_rsp_payload_data[31])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[30]  ( .D(
        iBusWishbone_DAT_MISO[30]), .CP(n7252), .Q(iBus_rsp_payload_data[30])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[29]  ( .D(
        iBusWishbone_DAT_MISO[29]), .CP(n7252), .Q(iBus_rsp_payload_data[29])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[28]  ( .D(
        iBusWishbone_DAT_MISO[28]), .CP(n7222), .Q(iBus_rsp_payload_data[28])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[27]  ( .D(
        iBusWishbone_DAT_MISO[27]), .CP(n7231), .Q(iBus_rsp_payload_data[27])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[26]  ( .D(
        iBusWishbone_DAT_MISO[26]), .CP(n7223), .Q(iBus_rsp_payload_data[26])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[25]  ( .D(
        iBusWishbone_DAT_MISO[25]), .CP(n7227), .Q(iBus_rsp_payload_data[25])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[24]  ( .D(
        iBusWishbone_DAT_MISO[24]), .CP(n7228), .Q(iBus_rsp_payload_data[24])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[23]  ( .D(
        iBusWishbone_DAT_MISO[23]), .CP(n7252), .Q(iBus_rsp_payload_data[23])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[22]  ( .D(
        iBusWishbone_DAT_MISO[22]), .CP(n7223), .Q(iBus_rsp_payload_data[22])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[21]  ( .D(
        iBusWishbone_DAT_MISO[21]), .CP(n7231), .Q(iBus_rsp_payload_data[21])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[20]  ( .D(
        iBusWishbone_DAT_MISO[20]), .CP(n7226), .Q(iBus_rsp_payload_data[20])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[19]  ( .D(
        iBusWishbone_DAT_MISO[19]), .CP(n7252), .Q(iBus_rsp_payload_data[19])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[18]  ( .D(
        iBusWishbone_DAT_MISO[18]), .CP(n7222), .Q(iBus_rsp_payload_data[18])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[17]  ( .D(
        iBusWishbone_DAT_MISO[17]), .CP(n7252), .Q(iBus_rsp_payload_data[17])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[16]  ( .D(
        iBusWishbone_DAT_MISO[16]), .CP(n7229), .Q(iBus_rsp_payload_data[16])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[15]  ( .D(
        iBusWishbone_DAT_MISO[15]), .CP(n7229), .Q(iBus_rsp_payload_data[15])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[14]  ( .D(
        iBusWishbone_DAT_MISO[14]), .CP(n7224), .Q(iBus_rsp_payload_data[14])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[13]  ( .D(
        iBusWishbone_DAT_MISO[13]), .CP(n7252), .Q(iBus_rsp_payload_data[13])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[12]  ( .D(
        iBusWishbone_DAT_MISO[12]), .CP(n7228), .Q(iBus_rsp_payload_data[12])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[11]  ( .D(
        iBusWishbone_DAT_MISO[11]), .CP(n7252), .Q(iBus_rsp_payload_data[11])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[10]  ( .D(
        iBusWishbone_DAT_MISO[10]), .CP(n7252), .Q(iBus_rsp_payload_data[10])
         );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[9]  ( .D(iBusWishbone_DAT_MISO[9]), 
        .CP(n7223), .Q(iBus_rsp_payload_data[9]) );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[8]  ( .D(iBusWishbone_DAT_MISO[8]), 
        .CP(n7227), .Q(iBus_rsp_payload_data[8]) );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[7]  ( .D(iBusWishbone_DAT_MISO[7]), 
        .CP(n7223), .Q(iBus_rsp_payload_data[7]) );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[6]  ( .D(iBusWishbone_DAT_MISO[6]), 
        .CP(n7226), .Q(iBus_rsp_payload_data[6]) );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[5]  ( .D(iBusWishbone_DAT_MISO[5]), 
        .CP(n7227), .Q(iBus_rsp_payload_data[5]) );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[4]  ( .D(iBusWishbone_DAT_MISO[4]), 
        .CP(n7223), .Q(iBus_rsp_payload_data[4]) );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[3]  ( .D(iBusWishbone_DAT_MISO[3]), 
        .CP(n7252), .Q(iBus_rsp_payload_data[3]) );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[2]  ( .D(iBusWishbone_DAT_MISO[2]), 
        .CP(n7252), .Q(iBus_rsp_payload_data[2]) );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[1]  ( .D(iBusWishbone_DAT_MISO[1]), 
        .CP(n7223), .Q(iBus_rsp_payload_data[1]) );
  dfnrq1 \iBusWishbone_DAT_MISO_regNext_reg[0]  ( .D(iBusWishbone_DAT_MISO[0]), 
        .CP(n7227), .Q(iBus_rsp_payload_data[0]) );
  dfnrq1 DebugPlugin_resetIt_reg ( .D(n4068), .CP(n7229), .Q(
        DebugPlugin_resetIt) );
  dfnrq1 DebugPlugin_resetIt_regNext_reg ( .D(DebugPlugin_resetIt), .CP(n7229), 
        .Q(debug_resetOut) );
  dfnrq1 DebugPlugin_debugUsed_reg ( .D(n6078), .CP(n7229), .Q(
        DebugPlugin_debugUsed) );
  dfnrq1 DebugPlugin_disableEbreak_reg ( .D(n6079), .CP(n7229), .Q(
        DebugPlugin_disableEbreak) );
  dfnrq1 DebugPlugin_stepIt_reg ( .D(n6075), .CP(n7229), .Q(DebugPlugin_stepIt) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][31]  ( .D(n6246), .CP(n7229), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[31]  ( .D(
        n6214), .CP(n7229), .Q(_zz_decode_LEGAL_INSTRUCTION_13_31) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[11]  ( .D(n5930), .CP(n7228), .Q(memory_REGFILE_WRITE_DATA[11]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[11]  ( .D(
        memory_REGFILE_WRITE_DATA[11]), .CP(n7228), .Q(
        writeBack_REGFILE_WRITE_DATA[11]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[10]  ( .D(n5929), .CP(n7228), .Q(memory_REGFILE_WRITE_DATA[10]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[10]  ( .D(
        memory_REGFILE_WRITE_DATA[10]), .CP(n7228), .Q(
        writeBack_REGFILE_WRITE_DATA[10]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[9]  ( .D(n5928), .CP(n7228), 
        .Q(memory_REGFILE_WRITE_DATA[9]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[9]  ( .D(
        memory_REGFILE_WRITE_DATA[9]), .CP(n7228), .Q(
        writeBack_REGFILE_WRITE_DATA[9]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[8]  ( .D(n5927), .CP(n7228), 
        .Q(memory_REGFILE_WRITE_DATA[8]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[8]  ( .D(
        memory_REGFILE_WRITE_DATA[8]), .CP(n7225), .Q(
        writeBack_REGFILE_WRITE_DATA[8]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[7]  ( .D(n5926), .CP(n7230), 
        .Q(memory_REGFILE_WRITE_DATA[7]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[7]  ( .D(
        memory_REGFILE_WRITE_DATA[7]), .CP(n7225), .Q(
        writeBack_REGFILE_WRITE_DATA[7]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[6]  ( .D(n5925), .CP(n7230), 
        .Q(memory_REGFILE_WRITE_DATA[6]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[6]  ( .D(
        memory_REGFILE_WRITE_DATA[6]), .CP(n7225), .Q(
        writeBack_REGFILE_WRITE_DATA[6]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[5]  ( .D(n5924), .CP(n7230), 
        .Q(memory_REGFILE_WRITE_DATA[5]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[5]  ( .D(
        memory_REGFILE_WRITE_DATA[5]), .CP(n7225), .Q(
        writeBack_REGFILE_WRITE_DATA[5]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[4]  ( .D(n5923), .CP(n7230), 
        .Q(memory_REGFILE_WRITE_DATA[4]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[4]  ( .D(
        memory_REGFILE_WRITE_DATA[4]), .CP(n7226), .Q(
        writeBack_REGFILE_WRITE_DATA[4]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[3]  ( .D(n5922), .CP(n7222), 
        .Q(memory_REGFILE_WRITE_DATA[3]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[3]  ( .D(
        memory_REGFILE_WRITE_DATA[3]), .CP(n7252), .Q(
        writeBack_REGFILE_WRITE_DATA[3]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[2]  ( .D(n5921), .CP(n7224), 
        .Q(memory_REGFILE_WRITE_DATA[2]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[2]  ( .D(
        memory_REGFILE_WRITE_DATA[2]), .CP(n7222), .Q(
        writeBack_REGFILE_WRITE_DATA[2]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[1]  ( .D(n5920), .CP(n7252), 
        .Q(memory_REGFILE_WRITE_DATA[1]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[1]  ( .D(
        memory_REGFILE_WRITE_DATA[1]), .CP(n7224), .Q(
        writeBack_REGFILE_WRITE_DATA[1]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[0]  ( .D(n5950), .CP(n7222), 
        .Q(memory_REGFILE_WRITE_DATA[0]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[0]  ( .D(
        memory_REGFILE_WRITE_DATA[0]), .CP(n7226), .Q(
        writeBack_REGFILE_WRITE_DATA[0]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[0]  ( .D(
        n6207), .CP(n7227), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[0]) );
  dfnrq1 \CsrPlugin_mtval_reg[0]  ( .D(n6039), .CP(n7222), .Q(
        CsrPlugin_mtval[0]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[0]  ( .D(n6165), .CP(n7231), .Q(_zz_CsrPlugin_csrMapping_readDataInit[0]) );
  dfnrq1 CsrPlugin_mip_MEIP_reg ( .D(N2210), .CP(n7229), .Q(CsrPlugin_mip_MEIP) );
  dfnrq1 \CsrPlugin_interrupt_code_reg[3]  ( .D(n4078), .CP(n7224), .Q(
        \CsrPlugin_interrupt_code[3] ) );
  dfnrq1 \CsrPlugin_mcause_exceptionCode_reg[3]  ( .D(n4074), .CP(n7222), .Q(
        CsrPlugin_mcause_exceptionCode[3]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[1]  ( .D(n4140), .CP(n7228), .Q(
        CsrPlugin_mtvec_base[1]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[3]  ( .D(n6116), .CP(n7228), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[3]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[3]  ( 
        .D(n5234), .CP(n7223), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[3]) );
  dfnrq1 \decode_to_execute_PC_reg[3]  ( .D(n5233), .CP(n7228), .Q(
        execute_PC[3]) );
  dfnrq1 \execute_LightShifterPlugin_amplitudeReg_reg[0]  ( .D(n4073), .CP(
        n7222), .Q(execute_LightShifterPlugin_amplitudeReg[0]) );
  dfnrq1 \execute_LightShifterPlugin_amplitudeReg_reg[1]  ( .D(n4072), .CP(
        n7223), .Q(execute_LightShifterPlugin_amplitudeReg[1]) );
  dfnrq1 \execute_LightShifterPlugin_amplitudeReg_reg[2]  ( .D(n4071), .CP(
        n7252), .Q(execute_LightShifterPlugin_amplitudeReg[2]) );
  dfnrq1 \execute_LightShifterPlugin_amplitudeReg_reg[3]  ( .D(n4070), .CP(
        n7224), .Q(execute_LightShifterPlugin_amplitudeReg[3]) );
  dfnrq1 \execute_LightShifterPlugin_amplitudeReg_reg[4]  ( .D(n4069), .CP(
        n7222), .Q(execute_LightShifterPlugin_amplitudeReg[4]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[29]  ( .D(n4112), .CP(n7227), .Q(
        CsrPlugin_mtvec_base[29]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[31]  ( .D(n6088), .CP(n7227), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[31]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[31]  ( 
        .D(n5318), .CP(n7227), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[31]) );
  dfnrq1 \decode_to_execute_PC_reg[31]  ( .D(n5317), .CP(n7227), .Q(
        execute_PC[31]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[30]  ( .D(n6089), .CP(n7227), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[30]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[30]  ( 
        .D(n5315), .CP(n7227), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[30]) );
  dfnrq1 \decode_to_execute_PC_reg[30]  ( .D(n5314), .CP(n7227), .Q(
        execute_PC[30]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[30]  ( .D(n5949), .CP(n7227), .Q(memory_REGFILE_WRITE_DATA[30]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[30]  ( .D(
        memory_REGFILE_WRITE_DATA[30]), .CP(n7227), .Q(
        writeBack_REGFILE_WRITE_DATA[30]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[29]  ( .D(n5948), .CP(n7227), .Q(memory_REGFILE_WRITE_DATA[29]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[29]  ( .D(
        memory_REGFILE_WRITE_DATA[29]), .CP(n7227), .Q(
        writeBack_REGFILE_WRITE_DATA[29]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[28]  ( .D(n5947), .CP(n7223), .Q(memory_REGFILE_WRITE_DATA[28]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[28]  ( .D(
        memory_REGFILE_WRITE_DATA[28]), .CP(n7227), .Q(
        writeBack_REGFILE_WRITE_DATA[28]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[27]  ( .D(n5946), .CP(n7223), .Q(memory_REGFILE_WRITE_DATA[27]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[27]  ( .D(
        memory_REGFILE_WRITE_DATA[27]), .CP(n7227), .Q(
        writeBack_REGFILE_WRITE_DATA[27]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[26]  ( .D(n5945), .CP(n7223), .Q(memory_REGFILE_WRITE_DATA[26]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[26]  ( .D(
        memory_REGFILE_WRITE_DATA[26]), .CP(n7223), .Q(
        writeBack_REGFILE_WRITE_DATA[26]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[25]  ( .D(n5944), .CP(n7223), .Q(memory_REGFILE_WRITE_DATA[25]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[25]  ( .D(
        memory_REGFILE_WRITE_DATA[25]), .CP(n7223), .Q(
        writeBack_REGFILE_WRITE_DATA[25]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[24]  ( .D(n5943), .CP(n7223), .Q(memory_REGFILE_WRITE_DATA[24]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[24]  ( .D(
        memory_REGFILE_WRITE_DATA[24]), .CP(n7223), .Q(
        writeBack_REGFILE_WRITE_DATA[24]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[23]  ( .D(n5942), .CP(n7223), .Q(memory_REGFILE_WRITE_DATA[23]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[23]  ( .D(
        memory_REGFILE_WRITE_DATA[23]), .CP(n7223), .Q(
        writeBack_REGFILE_WRITE_DATA[23]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[22]  ( .D(n5941), .CP(n7223), .Q(memory_REGFILE_WRITE_DATA[22]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[22]  ( .D(
        memory_REGFILE_WRITE_DATA[22]), .CP(n7226), .Q(
        writeBack_REGFILE_WRITE_DATA[22]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[21]  ( .D(n5940), .CP(n7226), .Q(memory_REGFILE_WRITE_DATA[21]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[21]  ( .D(
        memory_REGFILE_WRITE_DATA[21]), .CP(n7226), .Q(
        writeBack_REGFILE_WRITE_DATA[21]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[20]  ( .D(n5939), .CP(n7226), .Q(memory_REGFILE_WRITE_DATA[20]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[20]  ( .D(
        memory_REGFILE_WRITE_DATA[20]), .CP(n7226), .Q(
        writeBack_REGFILE_WRITE_DATA[20]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[19]  ( .D(n5938), .CP(n7226), .Q(memory_REGFILE_WRITE_DATA[19]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[19]  ( .D(
        memory_REGFILE_WRITE_DATA[19]), .CP(n7226), .Q(
        writeBack_REGFILE_WRITE_DATA[19]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[18]  ( .D(n5937), .CP(n7226), .Q(memory_REGFILE_WRITE_DATA[18]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[18]  ( .D(
        memory_REGFILE_WRITE_DATA[18]), .CP(n7225), .Q(
        writeBack_REGFILE_WRITE_DATA[18]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[17]  ( .D(n5936), .CP(n7225), .Q(memory_REGFILE_WRITE_DATA[17]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[17]  ( .D(
        memory_REGFILE_WRITE_DATA[17]), .CP(n7225), .Q(
        writeBack_REGFILE_WRITE_DATA[17]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[16]  ( .D(n5935), .CP(n7225), .Q(memory_REGFILE_WRITE_DATA[16]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[16]  ( .D(
        memory_REGFILE_WRITE_DATA[16]), .CP(n7225), .Q(
        writeBack_REGFILE_WRITE_DATA[16]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[15]  ( .D(n5934), .CP(n7225), .Q(memory_REGFILE_WRITE_DATA[15]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[15]  ( .D(
        memory_REGFILE_WRITE_DATA[15]), .CP(n7225), .Q(
        writeBack_REGFILE_WRITE_DATA[15]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[14]  ( .D(n5933), .CP(n7225), .Q(memory_REGFILE_WRITE_DATA[14]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[14]  ( .D(
        memory_REGFILE_WRITE_DATA[14]), .CP(n7224), .Q(
        writeBack_REGFILE_WRITE_DATA[14]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[13]  ( .D(n5932), .CP(n7224), .Q(memory_REGFILE_WRITE_DATA[13]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[13]  ( .D(
        memory_REGFILE_WRITE_DATA[13]), .CP(n7224), .Q(
        writeBack_REGFILE_WRITE_DATA[13]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[12]  ( .D(n5931), .CP(n7224), .Q(memory_REGFILE_WRITE_DATA[12]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[12]  ( .D(
        memory_REGFILE_WRITE_DATA[12]), .CP(n7224), .Q(
        writeBack_REGFILE_WRITE_DATA[12]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[12]  ( .D(
        n6187), .CP(n7224), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[12]) );
  dfnrq1 \CsrPlugin_mtval_reg[12]  ( .D(n6019), .CP(n7224), .Q(
        CsrPlugin_mtval[12]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[10]  ( .D(n4131), .CP(n7224), .Q(
        CsrPlugin_mtvec_base[10]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[12]  ( .D(n6107), .CP(n7226), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[12]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[2]  ( 
        .D(n5231), .CP(n7230), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[2]) );
  dfnrq1 \decode_to_execute_PC_reg[2]  ( .D(n5230), .CP(n7231), .Q(
        execute_PC[2]) );
  dfnrq1 \memory_to_writeBack_PC_reg[2]  ( .D(n5229), .CP(n7230), .Q(
        writeBack_PC[2]) );
  dfnrq1 \CsrPlugin_mepc_reg[2]  ( .D(n4109), .CP(n7230), .Q(CsrPlugin_mepc[2]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[0]  ( .D(
        n6245), .CP(n7225), .Q(_zz_decode_LEGAL_INSTRUCTION_1[0]) );
  dfnrq1 _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2_reg ( .D(n6119), 
        .CP(n7231), .Q(_zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1)
         );
  dfnrq1 DebugPlugin_haltIt_reg ( .D(n6074), .CP(n7230), .Q(DebugPlugin_haltIt) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[2]  ( .D(
        n6243), .CP(n7230), .Q(_zz_decode_LEGAL_INSTRUCTION_1[2]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[2]  ( .D(n5917), .CP(n7231), .Q(
        execute_INSTRUCTION[2]) );
  dfnrq1 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode_reg ( .D(N1781), .CP(n7230), .Q(CsrPlugin_exceptionPendings_0) );
  dfnrq1 \switch_Fetcher_l362_reg[1]  ( .D(n6169), .CP(n7230), .Q(
        switch_Fetcher_l362[1]) );
  dfnrq1 \switch_Fetcher_l362_reg[2]  ( .D(n6170), .CP(n7229), .Q(
        switch_Fetcher_l362[2]) );
  dfnrq1 \switch_Fetcher_l362_reg[0]  ( .D(n6171), .CP(n7231), .Q(
        switch_Fetcher_l362[0]) );
  dfnrq1 execute_arbitration_isValid_reg ( .D(n6166), .CP(n7224), .Q(
        execute_arbitration_isValid) );
  dfnrq1 memory_arbitration_isValid_reg ( .D(n6167), .CP(n7230), .Q(
        memory_arbitration_isValid) );
  dfnrq1 _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid_reg ( .D(
        n6120), .CP(n7230), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid) );
  dfnrq1 DebugPlugin_isPipBusy_reg ( .D(N2076), .CP(n7225), .Q(
        DebugPlugin_isPipBusy) );
  dfnrq1 DebugPlugin_godmode_reg ( .D(n6076), .CP(n7226), .Q(
        DebugPlugin_godmode) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_valid_reg  ( .D(n6080), .CP(n7230), 
        .Q(\IBusCachedPlugin_cache/lineLoader_valid ) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_cmdSent_reg  ( .D(n6082), .CP(
        n7228), .Q(\IBusCachedPlugin_cache/lineLoader_cmdSent ) );
  dfnrq1 \_zz_iBusWishbone_ADR_reg[0]  ( .D(n6174), .CP(n7230), .Q(
        iBusWishbone_ADR[0]) );
  dfnrq1 _zz_iBus_rsp_valid_reg ( .D(N1840), .CP(n7224), .Q(iBus_rsp_valid) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_wordIndex_reg[0]  ( .D(n6085), 
        .CP(n7225), .Q(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[0] )
         );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_wordIndex_reg[1]  ( .D(n6084), 
        .CP(n7228), .Q(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[1] )
         );
  dfnrq1 \_zz_iBusWishbone_ADR_reg[1]  ( .D(n6172), .CP(n7229), .Q(
        iBusWishbone_ADR[1]) );
  dfnrq1 \_zz_iBusWishbone_ADR_reg[2]  ( .D(n6173), .CP(n7226), .Q(
        iBusWishbone_ADR[2]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[31]  ( .D(n5915), .CP(
        n7225), .Q(iBusWishbone_ADR[29]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[30]  ( .D(n5914), .CP(
        n7228), .Q(iBusWishbone_ADR[28]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[12]  ( .D(n5896), .CP(
        n7229), .Q(iBusWishbone_ADR[10]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[5]  ( .D(n5889), .CP(
        n7231), .Q(iBusWishbone_ADR[3]) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][0]  ( .D(n5834), .CP(n7231), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][31]  ( .D(n5833), .CP(n7231), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][30]  ( .D(n5832), .CP(n7228), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][29]  ( .D(n5831), .CP(n7230), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][28]  ( .D(n5830), .CP(n7228), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][27]  ( .D(n5829), .CP(n7229), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][26]  ( .D(n5828), .CP(n7231), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][25]  ( .D(n5827), .CP(n7231), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][24]  ( .D(n5826), .CP(n7231), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][23]  ( .D(n5825), .CP(n7229), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][22]  ( .D(n5824), .CP(n7225), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][21]  ( .D(n5823), .CP(n7228), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][20]  ( .D(n5822), .CP(n7229), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][19]  ( .D(n5821), .CP(n7226), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][18]  ( .D(n5820), .CP(n7225), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][17]  ( .D(n5819), .CP(n7223), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][16]  ( .D(n5818), .CP(n7223), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][15]  ( .D(n5817), .CP(n7223), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][14]  ( .D(n5816), .CP(n7223), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][13]  ( .D(n5815), .CP(n7223), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][12]  ( .D(n5814), .CP(n7223), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][11]  ( .D(n5813), .CP(n7223), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][10]  ( .D(n5812), .CP(n7223), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][9]  ( .D(n5811), .CP(n7222), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][8]  ( .D(n5810), .CP(n7222), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][7]  ( .D(n5809), .CP(n7222), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][6]  ( .D(n5808), .CP(n7222), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][5]  ( .D(n5807), .CP(n7222), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][4]  ( .D(n5806), .CP(n7222), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][3]  ( .D(n5805), .CP(n7222), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][2]  ( .D(n5804), .CP(n7222), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[15][1]  ( .D(n5803), .CP(n7227), 
        .Q(\IBusCachedPlugin_cache/banks_0[15][1] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][0]  ( .D(n5770), .CP(n7223), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][31]  ( .D(n5769), .CP(n7231), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][30]  ( .D(n5768), .CP(n7252), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][29]  ( .D(n5767), .CP(n7229), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][28]  ( .D(n5766), .CP(n7226), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][27]  ( .D(n5765), .CP(n7252), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][26]  ( .D(n5764), .CP(n7224), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][25]  ( .D(n5763), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][24]  ( .D(n5762), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][23]  ( .D(n5761), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][22]  ( .D(n5760), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][21]  ( .D(n5759), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][20]  ( .D(n5758), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][19]  ( .D(n5757), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][18]  ( .D(n5756), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][17]  ( .D(n5755), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][16]  ( .D(n5754), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][15]  ( .D(n5753), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][14]  ( .D(n5752), .CP(clk), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][13]  ( .D(n5751), .CP(clk), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][12]  ( .D(n5750), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][11]  ( .D(n5749), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][10]  ( .D(n5748), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][9]  ( .D(n5747), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][8]  ( .D(n5746), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][7]  ( .D(n5745), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][6]  ( .D(n5744), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][5]  ( .D(n5743), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][4]  ( .D(n5742), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][3]  ( .D(n5741), .CP(clk), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][2]  ( .D(n5740), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[13][1]  ( .D(n5739), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[13][1] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][0]  ( .D(n5706), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][31]  ( .D(n5705), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][30]  ( .D(n5704), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][29]  ( .D(n5703), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][28]  ( .D(n5702), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][27]  ( .D(n5701), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][26]  ( .D(n5700), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][25]  ( .D(n5699), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][24]  ( .D(n5698), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][23]  ( .D(n5697), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][22]  ( .D(n5696), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][21]  ( .D(n5695), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][20]  ( .D(n5694), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][19]  ( .D(n5693), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][18]  ( .D(n5692), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][17]  ( .D(n5691), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][16]  ( .D(n5690), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][15]  ( .D(n5689), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][14]  ( .D(n5688), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][13]  ( .D(n5687), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][12]  ( .D(n5686), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][11]  ( .D(n5685), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][10]  ( .D(n5684), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][9]  ( .D(n5683), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][8]  ( .D(n5682), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][7]  ( .D(n5681), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][6]  ( .D(n5680), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][5]  ( .D(n5679), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][4]  ( .D(n5678), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][3]  ( .D(n5677), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][2]  ( .D(n5676), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[11][1]  ( .D(n5675), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[11][1] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][0]  ( .D(n5642), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][31]  ( .D(n5641), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][30]  ( .D(n5640), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][29]  ( .D(n5639), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][28]  ( .D(n5638), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][27]  ( .D(n5637), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][26]  ( .D(n5636), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][25]  ( .D(n5635), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][24]  ( .D(n5634), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][23]  ( .D(n5633), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][22]  ( .D(n5632), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][21]  ( .D(n5631), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][20]  ( .D(n5630), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][19]  ( .D(n5629), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][18]  ( .D(n5628), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][17]  ( .D(n5627), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][16]  ( .D(n5626), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][15]  ( .D(n5625), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][14]  ( .D(n5624), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][13]  ( .D(n5623), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][12]  ( .D(n5622), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][11]  ( .D(n5621), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][10]  ( .D(n5620), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][9]  ( .D(n5619), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][8]  ( .D(n5618), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][7]  ( .D(n5617), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][6]  ( .D(n5616), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][5]  ( .D(n5615), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][4]  ( .D(n5614), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][3]  ( .D(n5613), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][2]  ( .D(n5612), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[9][1]  ( .D(n5611), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[9][1] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][0]  ( .D(n5802), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][31]  ( .D(n5801), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][30]  ( .D(n5800), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][29]  ( .D(n5799), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][28]  ( .D(n5798), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][27]  ( .D(n5797), .CP(clk), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][26]  ( .D(n5796), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][25]  ( .D(n5795), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][24]  ( .D(n5794), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][23]  ( .D(n5793), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][22]  ( .D(n5792), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][21]  ( .D(n5791), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][20]  ( .D(n5790), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][19]  ( .D(n5789), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][18]  ( .D(n5788), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][17]  ( .D(n5787), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][16]  ( .D(n5786), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][15]  ( .D(n5785), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][14]  ( .D(n5784), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][13]  ( .D(n5783), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][12]  ( .D(n5782), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][11]  ( .D(n5781), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][10]  ( .D(n5780), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][9]  ( .D(n5779), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][8]  ( .D(n5778), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][7]  ( .D(n5777), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][6]  ( .D(n5776), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][5]  ( .D(n5775), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][4]  ( .D(n5774), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][3]  ( .D(n5773), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][2]  ( .D(n5772), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[14][1]  ( .D(n5771), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[14][1] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][0]  ( .D(n5738), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][31]  ( .D(n5737), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][30]  ( .D(n5736), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][29]  ( .D(n5735), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][28]  ( .D(n5734), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][27]  ( .D(n5733), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][26]  ( .D(n5732), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][25]  ( .D(n5731), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][24]  ( .D(n5730), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][23]  ( .D(n5729), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][22]  ( .D(n5728), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][21]  ( .D(n5727), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][20]  ( .D(n5726), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][19]  ( .D(n5725), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][18]  ( .D(n5724), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][17]  ( .D(n5723), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][16]  ( .D(n5722), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][15]  ( .D(n5721), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][14]  ( .D(n5720), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][13]  ( .D(n5719), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][12]  ( .D(n5718), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][11]  ( .D(n5717), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][10]  ( .D(n5716), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][9]  ( .D(n5715), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][8]  ( .D(n5714), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][7]  ( .D(n5713), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][6]  ( .D(n5712), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][5]  ( .D(n5711), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][4]  ( .D(n5710), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][3]  ( .D(n5709), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][2]  ( .D(n5708), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[12][1]  ( .D(n5707), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[12][1] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][0]  ( .D(n5674), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][31]  ( .D(n5673), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][30]  ( .D(n5672), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][29]  ( .D(n5671), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][28]  ( .D(n5670), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][27]  ( .D(n5669), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][26]  ( .D(n5668), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][25]  ( .D(n5667), .CP(clk), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][24]  ( .D(n5666), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][23]  ( .D(n5665), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][22]  ( .D(n5664), .CP(n7221), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][21]  ( .D(n5663), .CP(n7232), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][20]  ( .D(n5662), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][19]  ( .D(n5661), .CP(n7233), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][18]  ( .D(n5660), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][17]  ( .D(n5659), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][16]  ( .D(n5658), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][15]  ( .D(n5657), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][14]  ( .D(n5656), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][13]  ( .D(n5655), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][12]  ( .D(n5654), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][11]  ( .D(n5653), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][10]  ( .D(n5652), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][9]  ( .D(n5651), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][8]  ( .D(n5650), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][7]  ( .D(n5649), .CP(n7220), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][6]  ( .D(n5648), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][5]  ( .D(n5647), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][4]  ( .D(n5646), .CP(n7218), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][3]  ( .D(n5645), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][2]  ( .D(n5644), .CP(n7219), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[10][1]  ( .D(n5643), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[10][1] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][0]  ( .D(n5610), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][31]  ( .D(n5609), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][30]  ( .D(n5608), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][29]  ( .D(n5607), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][28]  ( .D(n5606), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][27]  ( .D(n5605), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][26]  ( .D(n5604), .CP(n7215), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][25]  ( .D(n5603), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][24]  ( .D(n5602), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][23]  ( .D(n5601), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][22]  ( .D(n5600), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][21]  ( .D(n5599), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][20]  ( .D(n5598), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][19]  ( .D(n5597), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][18]  ( .D(n5596), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][17]  ( .D(n5595), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][16]  ( .D(n5594), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][15]  ( .D(n5593), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][14]  ( .D(n5592), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][13]  ( .D(n5591), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][12]  ( .D(n5590), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][11]  ( .D(n5589), .CP(n7216), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][10]  ( .D(n5588), .CP(n7217), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][9]  ( .D(n5587), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][8]  ( .D(n5586), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][7]  ( .D(n5585), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][6]  ( .D(n5584), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][5]  ( .D(n5583), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][4]  ( .D(n5582), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][3]  ( .D(n5581), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][2]  ( .D(n5580), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[8][1]  ( .D(n5579), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[8][1] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][0]  ( .D(n5578), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][31]  ( .D(n5577), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][30]  ( .D(n5576), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][29]  ( .D(n5575), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][28]  ( .D(n5574), .CP(clk), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][27]  ( .D(n5573), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][26]  ( .D(n5572), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][25]  ( .D(n5571), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][24]  ( .D(n5570), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][23]  ( .D(n5569), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][22]  ( .D(n5568), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][21]  ( .D(n5567), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][20]  ( .D(n5566), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][19]  ( .D(n5565), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][18]  ( .D(n5564), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][17]  ( .D(n5563), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][16]  ( .D(n5562), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][15]  ( .D(n5561), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][14]  ( .D(n5560), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][13]  ( .D(n5559), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][12]  ( .D(n5558), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][11]  ( .D(n5557), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][10]  ( .D(n5556), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][9]  ( .D(n5555), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][8]  ( .D(n5554), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][7]  ( .D(n5553), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][6]  ( .D(n5552), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][5]  ( .D(n5551), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][4]  ( .D(n5550), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][3]  ( .D(n5549), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][2]  ( .D(n5548), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[7][1]  ( .D(n5547), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[7][1] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][0]  ( .D(n5514), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][31]  ( .D(n5513), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][30]  ( .D(n5512), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][29]  ( .D(n5511), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][28]  ( .D(n5510), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][27]  ( .D(n5509), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][26]  ( .D(n5508), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][25]  ( .D(n5507), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][24]  ( .D(n5506), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][23]  ( .D(n5505), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][22]  ( .D(n5504), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][21]  ( .D(n5503), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][20]  ( .D(n5502), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][19]  ( .D(n5501), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][18]  ( .D(n5500), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][17]  ( .D(n5499), .CP(n7146), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][16]  ( .D(n5498), .CP(n7164), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][15]  ( .D(n5497), .CP(n7191), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][14]  ( .D(n5496), .CP(n7200), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][13]  ( .D(n5495), .CP(n7137), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][12]  ( .D(n5494), .CP(n7182), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][11]  ( .D(n5493), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][10]  ( .D(n5492), .CP(n7123), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][9]  ( .D(n5491), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][8]  ( .D(n5490), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][7]  ( .D(n5489), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][6]  ( .D(n5488), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][5]  ( .D(n5487), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][4]  ( .D(n5486), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][3]  ( .D(n5485), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][2]  ( .D(n5484), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[5][1]  ( .D(n5483), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[5][1] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][0]  ( .D(n5450), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][31]  ( .D(n5449), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][30]  ( .D(n5448), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][29]  ( .D(n5447), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][28]  ( .D(n5446), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][27]  ( .D(n5445), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][26]  ( .D(n5444), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][25]  ( .D(n5443), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][24]  ( .D(n5442), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][23]  ( .D(n5441), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][22]  ( .D(n5440), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][21]  ( .D(n5439), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][20]  ( .D(n5438), .CP(n7213), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][19]  ( .D(n5437), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][18]  ( .D(n5436), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][17]  ( .D(n5435), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][16]  ( .D(n5434), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][15]  ( .D(n5433), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][14]  ( .D(n5432), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][13]  ( .D(n5431), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][12]  ( .D(n5430), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][11]  ( .D(n5429), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][10]  ( .D(n5428), .CP(n7214), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][9]  ( .D(n5427), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][8]  ( .D(n5426), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][7]  ( .D(n5425), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][6]  ( .D(n5424), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][5]  ( .D(n5423), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][4]  ( .D(n5422), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][3]  ( .D(n5421), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][2]  ( .D(n5420), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[3][1]  ( .D(n5419), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[3][1] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][0]  ( .D(n5386), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][31]  ( .D(n5385), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][30]  ( .D(n5384), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][29]  ( .D(n5383), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][28]  ( .D(n5382), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][27]  ( .D(n5381), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][26]  ( .D(n5380), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][25]  ( .D(n5379), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][24]  ( .D(n5378), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][23]  ( .D(n5377), .CP(n7155), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][22]  ( .D(n5376), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][21]  ( .D(n5375), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][20]  ( .D(n5374), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][19]  ( .D(n5373), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][18]  ( .D(n5372), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][17]  ( .D(n5371), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][16]  ( .D(n5370), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][15]  ( .D(n5369), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][14]  ( .D(n5368), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][13]  ( .D(n5367), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][12]  ( .D(n5366), .CP(n7173), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][11]  ( .D(n5365), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][10]  ( .D(n5364), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][9]  ( .D(n5363), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][8]  ( .D(n5362), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][7]  ( .D(n5361), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][6]  ( .D(n5360), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][5]  ( .D(n5359), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][4]  ( .D(n5358), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][3]  ( .D(n5357), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][2]  ( .D(n5356), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[1][1]  ( .D(n5355), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[1][1] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][0]  ( .D(n5546), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][31]  ( .D(n5545), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][30]  ( .D(n5544), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][29]  ( .D(n5543), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][28]  ( .D(n5542), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][27]  ( .D(n5541), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][26]  ( .D(n5540), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][25]  ( .D(n5539), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][24]  ( .D(n5538), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][23]  ( .D(n5537), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][22]  ( .D(n5536), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][21]  ( .D(n5535), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][20]  ( .D(n5534), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][19]  ( .D(n5533), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][18]  ( .D(n5532), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][17]  ( .D(n5531), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][16]  ( .D(n5530), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][15]  ( .D(n5529), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][14]  ( .D(n5528), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][13]  ( .D(n5527), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][12]  ( .D(n5526), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][11]  ( .D(n5525), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][10]  ( .D(n5524), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][9]  ( .D(n5523), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][8]  ( .D(n5522), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][7]  ( .D(n5521), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][6]  ( .D(n5520), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][5]  ( .D(n5519), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][4]  ( .D(n5518), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][3]  ( .D(n5517), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][2]  ( .D(n5516), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[6][1]  ( .D(n5515), .CP(n7234), 
        .Q(\IBusCachedPlugin_cache/banks_0[6][1] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][0]  ( .D(n5482), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][31]  ( .D(n5481), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][30]  ( .D(n5480), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][29]  ( .D(n5479), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][28]  ( .D(n5478), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][27]  ( .D(n5477), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][26]  ( .D(n5476), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][25]  ( .D(n5475), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][24]  ( .D(n5474), .CP(n7253), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][23]  ( .D(n5473), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][22]  ( .D(n5472), .CP(n7254), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][21]  ( .D(n5471), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][20]  ( .D(n5470), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][19]  ( .D(n5469), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][18]  ( .D(n5468), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][17]  ( .D(n5467), .CP(n7235), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][16]  ( .D(n5466), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][15]  ( .D(n5465), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][14]  ( .D(n5464), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][13]  ( .D(n5463), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][12]  ( .D(n5462), .CP(n7210), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][11]  ( .D(n5461), .CP(n7209), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][10]  ( .D(n5460), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][9]  ( .D(n5459), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][8]  ( .D(n5458), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][7]  ( .D(n5457), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][6]  ( .D(n5456), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][5]  ( .D(n5455), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][4]  ( .D(n5454), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][3]  ( .D(n5453), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][2]  ( .D(n5452), .CP(n7207), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[4][1]  ( .D(n5451), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[4][1] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][0]  ( .D(n5418), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][31]  ( .D(n5417), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][31] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][30]  ( .D(n5416), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][29]  ( .D(n5415), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][28]  ( .D(n5414), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][27]  ( .D(n5413), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][26]  ( .D(n5412), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][25]  ( .D(n5411), .CP(n7206), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][24]  ( .D(n5410), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][23]  ( .D(n5409), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][22]  ( .D(n5408), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][21]  ( .D(n5407), .CP(n7212), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][20]  ( .D(n5406), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][19]  ( .D(n5405), .CP(n7211), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][18]  ( .D(n5404), .CP(n7208), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][17]  ( .D(n5403), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][16]  ( .D(n5402), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][15]  ( .D(n5401), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][14]  ( .D(n5400), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][13]  ( .D(n5399), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][12]  ( .D(n5398), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][11]  ( .D(n5397), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][10]  ( .D(n5396), .CP(n7205), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][9]  ( .D(n5395), .CP(n7196), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][8]  ( .D(n5394), .CP(n7203), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][7]  ( .D(n5393), .CP(n7202), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][6]  ( .D(n5392), .CP(n7198), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][5]  ( .D(n5391), .CP(n7200), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][4]  ( .D(n5390), .CP(n7237), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][3]  ( .D(n5389), .CP(n7204), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][2]  ( .D(n5388), .CP(n7236), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[2][1]  ( .D(n5387), .CP(n7202), 
        .Q(\IBusCachedPlugin_cache/banks_0[2][1] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][0]  ( .D(n5354), .CP(n7203), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][30]  ( .D(n5353), .CP(n7255), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][30] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][29]  ( .D(n5352), .CP(n7236), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][29] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][28]  ( .D(n5351), .CP(n7201), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][28] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][27]  ( .D(n5350), .CP(n7201), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][26]  ( .D(n5349), .CP(n7197), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][25]  ( .D(n5348), .CP(n7196), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][24]  ( .D(n5347), .CP(n7255), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][23]  ( .D(n5346), .CP(n7203), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][22]  ( .D(n5345), .CP(n7202), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][21]  ( .D(n5344), .CP(n7255), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][20]  ( .D(n5343), .CP(n7203), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][19]  ( .D(n5342), .CP(n7255), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][18]  ( .D(n5341), .CP(n7236), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][17]  ( .D(n5340), .CP(n7201), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][16]  ( .D(n5339), .CP(n7201), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][15]  ( .D(n5338), .CP(n7197), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][14]  ( .D(n5337), .CP(n7236), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][13]  ( .D(n5336), .CP(n7200), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][12]  ( .D(n5335), .CP(n7196), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][11]  ( .D(n5334), .CP(n7255), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][10]  ( .D(n5333), .CP(n7197), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][9]  ( .D(n5332), .CP(n7199), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][8]  ( .D(n5331), .CP(n7236), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][7]  ( .D(n5330), .CP(n7236), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][6]  ( .D(n5329), .CP(n7236), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][5]  ( .D(n5328), .CP(n7236), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][4]  ( .D(n5327), .CP(n7199), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][3]  ( .D(n5326), .CP(n7203), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[3]  ( .D(
        n6242), .CP(n7236), .Q(_zz_decode_LEGAL_INSTRUCTION_1[3]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[3]  ( .D(n5918), .CP(n7196), .Q(
        execute_INSTRUCTION[3]) );
  dfnrq1 decode_to_execute_MEMORY_ENABLE_reg ( .D(n5981), .CP(n7236), .Q(
        execute_MEMORY_ENABLE) );
  dfnrq1 memory_to_writeBack_MEMORY_ENABLE_reg ( .D(memory_MEMORY_ENABLE), 
        .CP(n7236), .Q(writeBack_MEMORY_ENABLE) );
  dfnrq1 writeBack_arbitration_isValid_reg ( .D(n6168), .CP(n7199), .Q(
        lastStageIsValid) );
  dfnrq1 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack_reg ( .D(
        N1784), .CP(n7197), .Q(CsrPlugin_exceptionPendings_3) );
  dfnrq1 CsrPlugin_hadException_reg ( .D(N1792), .CP(n7236), .Q(
        CsrPlugin_hadException) );
  dfnrq1 CsrPlugin_mcause_interrupt_reg ( .D(n6040), .CP(n7199), .Q(
        CsrPlugin_mcause_interrupt) );
  dfnrq1 \memory_to_writeBack_PC_reg[31]  ( .D(n5316), .CP(n7197), .Q(
        writeBack_PC[31]) );
  dfnrq1 \memory_to_writeBack_PC_reg[30]  ( .D(n5313), .CP(n7196), .Q(
        writeBack_PC[30]) );
  dfnrq1 \memory_to_writeBack_PC_reg[5]  ( .D(n5238), .CP(n7204), .Q(
        writeBack_PC[5]) );
  dfnrq1 \CsrPlugin_mepc_reg[5]  ( .D(n4106), .CP(n7204), .Q(CsrPlugin_mepc[5]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[30]  ( .D(
        n6215), .CP(n7204), .Q(decode_INSTRUCTION_30) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[30]  ( .D(n5975), .CP(n7204), .Q(
        _zz__zz_execute_SRC2_3[10]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[29]  ( .D(
        n6216), .CP(n7204), .Q(_zz_decode_LEGAL_INSTRUCTION_13[29]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[29]  ( .D(n5974), .CP(n7204), .Q(
        _zz__zz_execute_SRC2_3[9]) );
  dfnrq1 \memory_to_writeBack_INSTRUCTION_reg[29]  ( .D(memory_INSTRUCTION_29), 
        .CP(n7204), .Q(_zz_lastStageRegFileWrite_payload_address_29) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[28]  ( .D(n5973), .CP(n7203), .Q(
        _zz__zz_execute_SRC2_3[8]) );
  dfnrq1 \memory_to_writeBack_INSTRUCTION_reg[28]  ( .D(memory_INSTRUCTION_28), 
        .CP(n7203), .Q(_zz_lastStageRegFileWrite_payload_address_28) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[27]  ( .D(
        n6218), .CP(n7203), .Q(_zz_decode_LEGAL_INSTRUCTION_13[27]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[27]  ( .D(n5972), .CP(n7203), .Q(
        _zz__zz_execute_SRC2_3[7]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[26]  ( .D(
        n6219), .CP(n7203), .Q(_zz_decode_LEGAL_INSTRUCTION_13[26]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[26]  ( .D(n5971), .CP(n7203), .Q(
        _zz__zz_execute_SRC2_3[6]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[25]  ( .D(
        n6220), .CP(n7203), .Q(_zz_decode_LEGAL_INSTRUCTION_13[25]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[25]  ( .D(n5970), .CP(n7203), .Q(
        _zz__zz_execute_SRC2_3[5]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[24]  ( .D(
        n6221), .CP(n7200), .Q(decode_INSTRUCTION_24) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[24]  ( .D(n5969), .CP(n7200), .Q(
        _zz__zz_execute_BranchPlugin_branch_src2_3) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[23]  ( .D(
        n6222), .CP(n7200), .Q(decode_INSTRUCTION_23) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[23]  ( .D(n5968), .CP(n7237), .Q(
        _zz__zz_execute_BranchPlugin_branch_src2_2) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[22]  ( .D(
        n6223), .CP(n7200), .Q(decode_INSTRUCTION_22) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[22]  ( .D(n5967), .CP(n7237), .Q(
        _zz__zz_execute_BranchPlugin_branch_src2_1) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[21]  ( .D(
        n6224), .CP(n7200), .Q(decode_INSTRUCTION_21) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[21]  ( .D(n5966), .CP(n7237), .Q(
        _zz__zz_execute_BranchPlugin_branch_src2_0) );
  dfnrq1 execute_CsrPlugin_csr_835_reg ( .D(n6005), .CP(n7198), .Q(
        execute_CsrPlugin_csr_835) );
  dfnrq1 \CsrPlugin_mepc_reg[0]  ( .D(n4111), .CP(n7204), .Q(CsrPlugin_mepc[0]) );
  dfnrq1 execute_CsrPlugin_csr_773_reg ( .D(n6002), .CP(n7198), .Q(
        execute_CsrPlugin_csr_773) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[20]  ( .D(n5965), .CP(n7204), .Q(
        _zz__zz_execute_BranchPlugin_branch_src2[10]) );
  dfnrq1 execute_CsrPlugin_csr_3008_reg ( .D(n6213), .CP(n7198), .Q(
        execute_CsrPlugin_csr_3008) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[12]  ( .D(n6145), .CP(
        n7204), .Q(_zz_CsrPlugin_csrMapping_readDataInit[12]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[3]  ( .D(n6136), .CP(n7255), .Q(_zz_CsrPlugin_csrMapping_readDataInit[3]) );
  dfnrq1 execute_CsrPlugin_csr_4032_reg ( .D(n6006), .CP(n7202), .Q(
        execute_CsrPlugin_csr_4032) );
  dfnrq1 execute_CsrPlugin_csr_834_reg ( .D(n6004), .CP(n7255), .Q(
        execute_CsrPlugin_csr_834) );
  dfnrq1 execute_CsrPlugin_csr_836_reg ( .D(n6000), .CP(n7237), .Q(
        execute_CsrPlugin_csr_836) );
  dfnrq1 CsrPlugin_mip_MSIP_reg ( .D(N2007), .CP(n7255), .Q(CsrPlugin_mip_MSIP) );
  dfnrq1 execute_CsrPlugin_csr_772_reg ( .D(n6001), .CP(n7255), .Q(
        execute_CsrPlugin_csr_772) );
  dfnrq1 CsrPlugin_mie_MSIE_reg ( .D(n6129), .CP(n7255), .Q(CsrPlugin_mie_MSIE) );
  dfnrq1 execute_CsrPlugin_csr_768_reg ( .D(n5999), .CP(n7204), .Q(
        execute_CsrPlugin_csr_768) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[19]  ( .D(
        n6226), .CP(n7255), .Q(decode_INSTRUCTION[19]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[19]  ( .D(n5964), .CP(n7255), .Q(
        _zz__zz_execute_SRC1_1[4]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[18]  ( .D(
        n6227), .CP(n7255), .Q(decode_INSTRUCTION[18]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[18]  ( .D(n5963), .CP(n7255), .Q(
        _zz__zz_execute_SRC1_1[3]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[17]  ( .D(
        n6228), .CP(n7200), .Q(decode_INSTRUCTION[17]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[17]  ( .D(n5962), .CP(n7237), .Q(
        _zz__zz_execute_SRC1_1[2]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[16]  ( .D(
        n6229), .CP(n7255), .Q(decode_INSTRUCTION[16]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[16]  ( .D(n5961), .CP(n7255), .Q(
        _zz__zz_execute_SRC1_1[1]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[15]  ( .D(
        n6230), .CP(n7237), .Q(decode_INSTRUCTION[15]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[15]  ( .D(n5960), .CP(n7201), .Q(
        _zz__zz_execute_SRC1_1[0]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[14]  ( .D(n5959), .CP(n7237), .Q(
        _zz__zz_execute_BranchPlugin_branch_src2[13]) );
  dfnrq1 \memory_to_writeBack_INSTRUCTION_reg[14]  ( .D(memory_INSTRUCTION[14]), .CP(n7201), .Q(_zz_lastStageRegFileWrite_payload_address[14]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[13]  ( .D(
        n6232), .CP(n7236), .Q(_zz_decode_LEGAL_INSTRUCTION_1_13) );
  dfnrq1 decode_to_execute_CSR_WRITE_OPCODE_reg ( .D(n5998), .CP(n7202), .Q(
        execute_CSR_WRITE_OPCODE) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[13]  ( .D(n5958), .CP(n7237), .Q(
        _zz__zz_execute_BranchPlugin_branch_src2[12]) );
  dfnrq1 \memory_to_writeBack_INSTRUCTION_reg[13]  ( .D(memory_INSTRUCTION[13]), .CP(n7237), .Q(_zz_lastStageRegFileWrite_payload_address[13]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[12]  ( .D(
        n6233), .CP(n7236), .Q(_zz_decode_LEGAL_INSTRUCTION_7_12) );
  dfnrq1 \decode_to_execute_ALU_BITWISE_CTRL_reg[1]  ( .D(n5988), .CP(n7204), 
        .Q(execute_ALU_BITWISE_CTRL[1]) );
  dfnrq1 \memory_to_writeBack_INSTRUCTION_reg[12]  ( .D(memory_INSTRUCTION[12]), .CP(n7197), .Q(_zz_lastStageRegFileWrite_payload_address[12]) );
  dfnrq1 \decode_to_execute_ALU_BITWISE_CTRL_reg[0]  ( .D(n5989), .CP(n7237), 
        .Q(execute_ALU_BITWISE_CTRL[0]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[11]  ( .D(
        n6234), .CP(n7236), .Q(decode_INSTRUCTION_11) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[11]  ( .D(n5957), .CP(n7237), .Q(
        _zz__zz_execute_SRC2_3[4]) );
  dfnrq1 \memory_to_writeBack_INSTRUCTION_reg[11]  ( .D(memory_INSTRUCTION[11]), .CP(n7196), .Q(_zz_lastStageRegFileWrite_payload_address[11]) );
  dfnrq1 \HazardSimplePlugin_writeBackBuffer_payload_address_reg[4]  ( .D(
        _zz_lastStageRegFileWrite_payload_address[11]), .CP(n7237), .Q(
        HazardSimplePlugin_writeBackBuffer_payload_address[4]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[10]  ( .D(
        n6235), .CP(n7198), .Q(decode_INSTRUCTION_10) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[10]  ( .D(n5956), .CP(n7200), .Q(
        _zz__zz_execute_SRC2_3[3]) );
  dfnrq1 \memory_to_writeBack_INSTRUCTION_reg[10]  ( .D(memory_INSTRUCTION[10]), .CP(n7203), .Q(_zz_lastStageRegFileWrite_payload_address[10]) );
  dfnrq1 \HazardSimplePlugin_writeBackBuffer_payload_address_reg[3]  ( .D(
        _zz_lastStageRegFileWrite_payload_address[10]), .CP(n7204), .Q(
        HazardSimplePlugin_writeBackBuffer_payload_address[3]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[9]  ( .D(
        n6236), .CP(n7198), .Q(decode_INSTRUCTION_9) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[9]  ( .D(n5955), .CP(n7200), .Q(
        _zz__zz_execute_SRC2_3[2]) );
  dfnrq1 \HazardSimplePlugin_writeBackBuffer_payload_address_reg[2]  ( .D(
        _zz_lastStageRegFileWrite_payload_address[9]), .CP(n7202), .Q(
        HazardSimplePlugin_writeBackBuffer_payload_address[2]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[8]  ( .D(
        n6237), .CP(n7202), .Q(decode_INSTRUCTION_8) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[8]  ( .D(n5954), .CP(n7202), .Q(
        _zz__zz_execute_SRC2_3[1]) );
  dfnrq1 \HazardSimplePlugin_writeBackBuffer_payload_address_reg[1]  ( .D(
        _zz_lastStageRegFileWrite_payload_address[8]), .CP(n7202), .Q(
        HazardSimplePlugin_writeBackBuffer_payload_address[1]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[7]  ( .D(
        n6238), .CP(n7202), .Q(decode_INSTRUCTION_7) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[7]  ( .D(n5953), .CP(n7202), .Q(
        _zz__zz_execute_SRC2_3[0]) );
  dfnrq1 \memory_to_writeBack_INSTRUCTION_reg[7]  ( .D(memory_INSTRUCTION[7]), 
        .CP(n7202), .Q(_zz_lastStageRegFileWrite_payload_address[7]) );
  dfnrq1 \HazardSimplePlugin_writeBackBuffer_payload_address_reg[0]  ( .D(
        _zz_lastStageRegFileWrite_payload_address[7]), .CP(n7201), .Q(
        HazardSimplePlugin_writeBackBuffer_payload_address[0]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[6]  ( .D(n5952), .CP(n7201), .Q(
        execute_INSTRUCTION[6]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[5]  ( .D(
        n6240), .CP(n7201), .Q(_zz_decode_LEGAL_INSTRUCTION_1[5]) );
  dfnrq1 \decode_to_execute_SRC2_CTRL_reg[0]  ( .D(n5985), .CP(n7201), .Q(
        execute_SRC2_CTRL[0]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[5]  ( .D(n5951), .CP(n7201), .Q(
        execute_INSTRUCTION[5]) );
  dfnrq1 decode_to_execute_SRC_USE_SUB_LESS_reg ( .D(n5980), .CP(n7201), .Q(
        execute_SRC_USE_SUB_LESS) );
  dfnrq1 \decode_to_execute_ENV_CTRL_reg[0]  ( .D(n5996), .CP(n7200), .Q(
        execute_ENV_CTRL[0]) );
  dfnrq1 \memory_to_writeBack_ENV_CTRL_reg[0]  ( .D(memory_ENV_CTRL[0]), .CP(
        n7200), .Q(writeBack_ENV_CTRL[0]) );
  dfnrq1 decode_to_execute_DO_EBREAK_reg ( .D(n6073), .CP(n7200), .Q(
        execute_DO_EBREAK) );
  dfnrq1 \decode_to_execute_ENV_CTRL_reg[1]  ( .D(n5995), .CP(n7200), .Q(
        execute_ENV_CTRL[1]) );
  dfnrq1 \memory_to_writeBack_ENV_CTRL_reg[1]  ( .D(memory_ENV_CTRL[1]), .CP(
        n7200), .Q(writeBack_ENV_CTRL[1]) );
  dfnrq1 \CsrPlugin_mstatus_MPP_reg[1]  ( .D(n6126), .CP(n7200), .Q(
        CsrPlugin_mstatus_MPP[1]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_code_reg[2]  ( .D(n6209), .CP(n7200), .Q(CsrPlugin_exceptionPortCtrl_exceptionContext_code[2]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_code_reg[0]  ( .D(n6211), .CP(n7200), .Q(CsrPlugin_exceptionPortCtrl_exceptionContext_code[0]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_code_reg[3]  ( .D(n6210), .CP(n7204), .Q(CsrPlugin_exceptionPortCtrl_exceptionContext_code[3]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_code_reg[1]  ( .D(n6208), .CP(n7197), .Q(CsrPlugin_exceptionPortCtrl_exceptionContext_code[1]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[30]  ( .D(
        n6205), .CP(n7201), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[30]) );
  dfnrq1 \CsrPlugin_mtval_reg[30]  ( .D(n6037), .CP(n7255), .Q(
        CsrPlugin_mtval[30]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[3]  ( .D(
        n6178), .CP(n7236), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[3]) );
  dfnrq1 \CsrPlugin_mtval_reg[3]  ( .D(n6010), .CP(n7203), .Q(
        CsrPlugin_mtval[3]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[2]  ( .D(
        n6177), .CP(n7202), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[2]) );
  dfnrq1 \CsrPlugin_mtval_reg[2]  ( .D(n6009), .CP(n7196), .Q(
        CsrPlugin_mtval[2]) );
  dfnrq1 execute_LightShifterPlugin_isActive_reg ( .D(n6123), .CP(n7199), .Q(
        execute_LightShifterPlugin_isActive) );
  dfnrq1 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute_reg ( .D(
        N1782), .CP(n7199), .Q(CsrPlugin_exceptionPendings_1) );
  dfnrq1 decode_to_execute_IS_CSR_reg ( .D(n5994), .CP(n7199), .Q(
        execute_IS_CSR) );
  dfnrq1 decode_to_execute_SRC2_FORCE_ZERO_reg ( .D(n5997), .CP(n7199), .Q(
        execute_SRC2_FORCE_ZERO) );
  dfnrq1 \decode_to_execute_SHIFT_CTRL_reg[0]  ( .D(n5991), .CP(n7199), .Q(
        execute_SHIFT_CTRL[0]) );
  dfnrq1 \decode_to_execute_SHIFT_CTRL_reg[1]  ( .D(n5990), .CP(n7199), .Q(
        execute_SHIFT_CTRL[1]) );
  dfnrq1 decode_to_execute_REGFILE_WRITE_VALID_reg ( .D(n5986), .CP(n7199), 
        .Q(execute_REGFILE_WRITE_VALID) );
  dfnrq1 memory_to_writeBack_REGFILE_WRITE_VALID_reg ( .D(
        memory_REGFILE_WRITE_VALID), .CP(n7199), .Q(
        writeBack_REGFILE_WRITE_VALID) );
  dfnrq1 HazardSimplePlugin_writeBackBuffer_valid_reg ( .D(N1771), .CP(n7236), 
        .Q(HazardSimplePlugin_writeBackBuffer_valid) );
  dfnrq1 \decode_to_execute_ALU_CTRL_reg[0]  ( .D(n5983), .CP(n7201), .Q(
        execute_ALU_CTRL[0]) );
  dfnrq1 \decode_to_execute_ALU_CTRL_reg[1]  ( .D(n5982), .CP(n7197), .Q(
        execute_ALU_CTRL[1]) );
  dfnrq1 \decode_to_execute_SRC1_CTRL_reg[0]  ( .D(n5979), .CP(n7197), .Q(
        execute_SRC1_CTRL[0]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[4]  ( .D(n5919), .CP(n7196), .Q(
        execute_INSTRUCTION[4]) );
  dfnrq1 \decode_to_execute_BRANCH_CTRL_reg[0]  ( .D(n5993), .CP(n7203), .Q(
        execute_BRANCH_CTRL[0]) );
  dfnrq1 decode_to_execute_SRC_LESS_UNSIGNED_reg ( .D(n5987), .CP(n7202), .Q(
        execute_SRC_LESS_UNSIGNED) );
  dfnrq1 \decode_to_execute_SRC2_CTRL_reg[1]  ( .D(n5984), .CP(n7198), .Q(
        execute_SRC2_CTRL[1]) );
  dfnrq1 \decode_to_execute_BRANCH_CTRL_reg[1]  ( .D(n5992), .CP(n7204), .Q(
        execute_BRANCH_CTRL[1]) );
  dfnrq1 \decode_to_execute_SRC1_CTRL_reg[1]  ( .D(n5978), .CP(n7201), .Q(
        execute_SRC1_CTRL[1]) );
  dfnrq1 \memory_to_writeBack_MEMORY_ADDRESS_LOW_reg[0]  ( .D(
        memory_MEMORY_ADDRESS_LOW[0]), .CP(n7255), .Q(
        writeBack_MEMORY_ADDRESS_LOW[0]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[1]  ( .D(n6071), .CP(n7197), .Q(
        DebugPlugin_busReadDataReg[1]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][1]  ( .D(n5197), .CP(n7196), .Q(
        \RegFilePlugin_regFile[31][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][1]  ( .D(n5165), .CP(n7203), .Q(
        \RegFilePlugin_regFile[30][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][1]  ( .D(n5133), .CP(n7202), .Q(
        \RegFilePlugin_regFile[29][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][1]  ( .D(n5101), .CP(n7198), .Q(
        \RegFilePlugin_regFile[28][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][1]  ( .D(n5069), .CP(n7199), .Q(
        \RegFilePlugin_regFile[27][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][1]  ( .D(n5037), .CP(n7202), .Q(
        \RegFilePlugin_regFile[26][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][1]  ( .D(n5005), .CP(n7203), .Q(
        \RegFilePlugin_regFile[25][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][1]  ( .D(n4973), .CP(n7196), .Q(
        \RegFilePlugin_regFile[24][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][1]  ( .D(n4941), .CP(n7197), .Q(
        \RegFilePlugin_regFile[23][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][1]  ( .D(n4909), .CP(n7201), .Q(
        \RegFilePlugin_regFile[22][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][1]  ( .D(n4877), .CP(n7237), .Q(
        \RegFilePlugin_regFile[21][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][1]  ( .D(n4845), .CP(n7202), .Q(
        \RegFilePlugin_regFile[20][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][1]  ( .D(n4813), .CP(n7198), .Q(
        \RegFilePlugin_regFile[19][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][1]  ( .D(n4781), .CP(n7198), .Q(
        \RegFilePlugin_regFile[18][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][1]  ( .D(n4749), .CP(n7198), .Q(
        \RegFilePlugin_regFile[17][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][1]  ( .D(n4717), .CP(n7198), .Q(
        \RegFilePlugin_regFile[16][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][1]  ( .D(n4685), .CP(n7198), .Q(
        \RegFilePlugin_regFile[15][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][1]  ( .D(n4653), .CP(n7198), .Q(
        \RegFilePlugin_regFile[14][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][1]  ( .D(n4621), .CP(n7198), .Q(
        \RegFilePlugin_regFile[13][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][1]  ( .D(n4589), .CP(n7198), .Q(
        \RegFilePlugin_regFile[12][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][1]  ( .D(n4557), .CP(n7197), .Q(
        \RegFilePlugin_regFile[11][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][1]  ( .D(n4525), .CP(n7197), .Q(
        \RegFilePlugin_regFile[10][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][1]  ( .D(n4493), .CP(n7197), .Q(
        \RegFilePlugin_regFile[9][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][1]  ( .D(n4461), .CP(n7197), .Q(
        \RegFilePlugin_regFile[8][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][1]  ( .D(n4429), .CP(n7197), .Q(
        \RegFilePlugin_regFile[7][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][1]  ( .D(n4397), .CP(n7197), .Q(
        \RegFilePlugin_regFile[6][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][1]  ( .D(n4365), .CP(n7197), .Q(
        \RegFilePlugin_regFile[5][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][1]  ( .D(n4333), .CP(n7197), .Q(
        \RegFilePlugin_regFile[4][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][1]  ( .D(n4301), .CP(n7196), .Q(
        \RegFilePlugin_regFile[3][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][1]  ( .D(n4269), .CP(n7199), .Q(
        \RegFilePlugin_regFile[2][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][1]  ( .D(n4237), .CP(n7203), .Q(
        \RegFilePlugin_regFile[1][1] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][1]  ( .D(n4144), .CP(n7199), .Q(
        \RegFilePlugin_regFile[0][1] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[1]  ( .D(N853), .CP(n7202), .Q(
        _zz_RegFilePlugin_regFile_port0[1]) );
  dfnrq1 \decode_to_execute_RS1_reg[1]  ( .D(n4143), .CP(n7199), .Q(
        execute_RS1[1]) );
  dfnrq1 \memory_to_writeBack_MEMORY_ADDRESS_LOW_reg[1]  ( .D(
        memory_MEMORY_ADDRESS_LOW[1]), .CP(n7198), .Q(
        writeBack_MEMORY_ADDRESS_LOW[1]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[0]  ( .D(n6072), .CP(n7199), .Q(
        DebugPlugin_busReadDataReg[0]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][0]  ( .D(n5228), .CP(n7196), .Q(
        \RegFilePlugin_regFile[31][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][0]  ( .D(n5196), .CP(n7196), .Q(
        \RegFilePlugin_regFile[30][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][0]  ( .D(n5164), .CP(n7196), .Q(
        \RegFilePlugin_regFile[29][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][0]  ( .D(n5132), .CP(n7196), .Q(
        \RegFilePlugin_regFile[28][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][0]  ( .D(n5100), .CP(n7196), .Q(
        \RegFilePlugin_regFile[27][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][0]  ( .D(n5068), .CP(n7196), .Q(
        \RegFilePlugin_regFile[26][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][0]  ( .D(n5036), .CP(n7196), .Q(
        \RegFilePlugin_regFile[25][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][0]  ( .D(n5004), .CP(n7196), .Q(
        \RegFilePlugin_regFile[24][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][0]  ( .D(n4972), .CP(n7187), .Q(
        \RegFilePlugin_regFile[23][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][0]  ( .D(n4940), .CP(n7194), .Q(
        \RegFilePlugin_regFile[22][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][0]  ( .D(n4908), .CP(n7193), .Q(
        \RegFilePlugin_regFile[21][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][0]  ( .D(n4876), .CP(n7189), .Q(
        \RegFilePlugin_regFile[20][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][0]  ( .D(n4844), .CP(n7191), .Q(
        \RegFilePlugin_regFile[19][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][0]  ( .D(n4812), .CP(n7239), .Q(
        \RegFilePlugin_regFile[18][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][0]  ( .D(n4780), .CP(n7195), .Q(
        \RegFilePlugin_regFile[17][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][0]  ( .D(n4748), .CP(n7238), .Q(
        \RegFilePlugin_regFile[16][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][0]  ( .D(n4716), .CP(n7193), .Q(
        \RegFilePlugin_regFile[15][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][0]  ( .D(n4684), .CP(n7194), .Q(
        \RegFilePlugin_regFile[14][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][0]  ( .D(n4652), .CP(n7256), .Q(
        \RegFilePlugin_regFile[13][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][0]  ( .D(n4620), .CP(n7238), .Q(
        \RegFilePlugin_regFile[12][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][0]  ( .D(n4588), .CP(n7192), .Q(
        \RegFilePlugin_regFile[11][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][0]  ( .D(n4556), .CP(n7192), .Q(
        \RegFilePlugin_regFile[10][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][0]  ( .D(n4524), .CP(n7188), .Q(
        \RegFilePlugin_regFile[9][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][0]  ( .D(n4492), .CP(n7187), .Q(
        \RegFilePlugin_regFile[8][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][0]  ( .D(n4460), .CP(n7256), .Q(
        \RegFilePlugin_regFile[7][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][0]  ( .D(n4428), .CP(n7194), .Q(
        \RegFilePlugin_regFile[6][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][0]  ( .D(n4396), .CP(n7193), .Q(
        \RegFilePlugin_regFile[5][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][0]  ( .D(n4364), .CP(n7256), .Q(
        \RegFilePlugin_regFile[4][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][0]  ( .D(n4332), .CP(n7194), .Q(
        \RegFilePlugin_regFile[3][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][0]  ( .D(n4300), .CP(n7256), .Q(
        \RegFilePlugin_regFile[2][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][0]  ( .D(n4268), .CP(n7238), .Q(
        \RegFilePlugin_regFile[1][0] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][0]  ( .D(n4236), .CP(n7192), .Q(
        \RegFilePlugin_regFile[0][0] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[0]  ( .D(N854), .CP(n7192), .Q(
        _zz_RegFilePlugin_regFile_port0[0]) );
  dfnrq1 \decode_to_execute_RS1_reg[0]  ( .D(n4235), .CP(n7188), .Q(
        execute_RS1[0]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[0]  ( .D(N887), .CP(n7238), .Q(
        _zz_RegFilePlugin_regFile_port1[0]) );
  dfnrq1 \decode_to_execute_RS2_reg[0]  ( .D(n6007), .CP(n7191), .Q(
        execute_RS2[0]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[30]  ( .D(n6042), .CP(n7187), .Q(
        debug_bus_rsp_data[30]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][30]  ( .D(n5226), .CP(n7256), .Q(
        \RegFilePlugin_regFile[31][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][30]  ( .D(n5194), .CP(n7188), .Q(
        \RegFilePlugin_regFile[30][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][30]  ( .D(n5162), .CP(n7190), .Q(
        \RegFilePlugin_regFile[29][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][30]  ( .D(n5130), .CP(n7238), .Q(
        \RegFilePlugin_regFile[28][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][30]  ( .D(n5098), .CP(n7238), .Q(
        \RegFilePlugin_regFile[27][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][30]  ( .D(n5066), .CP(n7238), .Q(
        \RegFilePlugin_regFile[26][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][30]  ( .D(n5034), .CP(n7238), .Q(
        \RegFilePlugin_regFile[25][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][30]  ( .D(n5002), .CP(n7190), .Q(
        \RegFilePlugin_regFile[24][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][30]  ( .D(n4970), .CP(n7194), .Q(
        \RegFilePlugin_regFile[23][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][30]  ( .D(n4938), .CP(n7238), .Q(
        \RegFilePlugin_regFile[22][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][30]  ( .D(n4906), .CP(n7187), .Q(
        \RegFilePlugin_regFile[21][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][30]  ( .D(n4874), .CP(n7238), .Q(
        \RegFilePlugin_regFile[20][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][30]  ( .D(n4842), .CP(n7238), .Q(
        \RegFilePlugin_regFile[19][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][30]  ( .D(n4810), .CP(n7190), .Q(
        \RegFilePlugin_regFile[18][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][30]  ( .D(n4778), .CP(n7188), .Q(
        \RegFilePlugin_regFile[17][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][30]  ( .D(n4746), .CP(n7238), .Q(
        \RegFilePlugin_regFile[16][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][30]  ( .D(n4714), .CP(n7190), .Q(
        \RegFilePlugin_regFile[15][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][30]  ( .D(n4682), .CP(n7188), .Q(
        \RegFilePlugin_regFile[14][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][30]  ( .D(n4650), .CP(n7187), .Q(
        \RegFilePlugin_regFile[13][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][30]  ( .D(n4618), .CP(n7195), .Q(
        \RegFilePlugin_regFile[12][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][30]  ( .D(n4586), .CP(n7195), .Q(
        \RegFilePlugin_regFile[11][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][30]  ( .D(n4554), .CP(n7195), .Q(
        \RegFilePlugin_regFile[10][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][30]  ( .D(n4522), .CP(n7195), .Q(
        \RegFilePlugin_regFile[9][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][30]  ( .D(n4490), .CP(n7195), .Q(
        \RegFilePlugin_regFile[8][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][30]  ( .D(n4458), .CP(n7195), .Q(
        \RegFilePlugin_regFile[7][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][30]  ( .D(n4426), .CP(n7195), .Q(
        \RegFilePlugin_regFile[6][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][30]  ( .D(n4394), .CP(n7195), .Q(
        \RegFilePlugin_regFile[5][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][30]  ( .D(n4362), .CP(n7194), .Q(
        \RegFilePlugin_regFile[4][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][30]  ( .D(n4330), .CP(n7194), .Q(
        \RegFilePlugin_regFile[3][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][30]  ( .D(n4298), .CP(n7194), .Q(
        \RegFilePlugin_regFile[2][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][30]  ( .D(n4266), .CP(n7194), .Q(
        \RegFilePlugin_regFile[1][30] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][30]  ( .D(n4231), .CP(n7194), .Q(
        \RegFilePlugin_regFile[0][30] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[30]  ( .D(N824), .CP(n7194), .Q(
        _zz_RegFilePlugin_regFile_port0[30]) );
  dfnrq1 \decode_to_execute_RS1_reg[30]  ( .D(n4230), .CP(n7194), .Q(
        execute_RS1[30]) );
  dfnrq1 \CsrPlugin_mepc_reg[30]  ( .D(n4081), .CP(n7194), .Q(
        CsrPlugin_mepc[30]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[30]  ( .D(n6163), .CP(
        n7191), .Q(_zz_CsrPlugin_csrMapping_readDataInit[30]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[28]  ( .D(n4113), .CP(n7191), .Q(
        CsrPlugin_mtvec_base[28]) );
  dfnrq1 \execute_to_memory_REGFILE_WRITE_DATA_reg[31]  ( .D(n6212), .CP(n7191), .Q(memory_REGFILE_WRITE_DATA[31]) );
  dfnrq1 \memory_to_writeBack_REGFILE_WRITE_DATA_reg[31]  ( .D(
        memory_REGFILE_WRITE_DATA[31]), .CP(n7239), .Q(
        writeBack_REGFILE_WRITE_DATA[31]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[31]  ( .D(n6041), .CP(n7191), .Q(
        debug_bus_rsp_data[31]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][31]  ( .D(n5227), .CP(n7239), .Q(
        \RegFilePlugin_regFile[31][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][31]  ( .D(n5195), .CP(n7191), .Q(
        \RegFilePlugin_regFile[30][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][31]  ( .D(n5163), .CP(n7239), .Q(
        \RegFilePlugin_regFile[29][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][31]  ( .D(n5131), .CP(n7189), .Q(
        \RegFilePlugin_regFile[28][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][31]  ( .D(n5099), .CP(n7189), .Q(
        \RegFilePlugin_regFile[27][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][31]  ( .D(n5067), .CP(n7189), .Q(
        \RegFilePlugin_regFile[26][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][31]  ( .D(n5035), .CP(n7195), .Q(
        \RegFilePlugin_regFile[25][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][31]  ( .D(n5003), .CP(n7189), .Q(
        \RegFilePlugin_regFile[24][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][31]  ( .D(n4971), .CP(n7195), .Q(
        \RegFilePlugin_regFile[23][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][31]  ( .D(n4939), .CP(n7189), .Q(
        \RegFilePlugin_regFile[22][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][31]  ( .D(n4907), .CP(n7195), .Q(
        \RegFilePlugin_regFile[21][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][31]  ( .D(n4875), .CP(n7256), .Q(
        \RegFilePlugin_regFile[20][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][31]  ( .D(n4843), .CP(n7193), .Q(
        \RegFilePlugin_regFile[19][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][31]  ( .D(n4811), .CP(n7256), .Q(
        \RegFilePlugin_regFile[18][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][31]  ( .D(n4779), .CP(n7239), .Q(
        \RegFilePlugin_regFile[17][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][31]  ( .D(n4747), .CP(n7256), .Q(
        \RegFilePlugin_regFile[16][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][31]  ( .D(n4715), .CP(n7256), .Q(
        \RegFilePlugin_regFile[15][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][31]  ( .D(n4683), .CP(n7256), .Q(
        \RegFilePlugin_regFile[14][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][31]  ( .D(n4651), .CP(n7195), .Q(
        \RegFilePlugin_regFile[13][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][31]  ( .D(n4619), .CP(n7256), .Q(
        \RegFilePlugin_regFile[12][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][31]  ( .D(n4587), .CP(n7256), .Q(
        \RegFilePlugin_regFile[11][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][31]  ( .D(n4555), .CP(n7256), .Q(
        \RegFilePlugin_regFile[10][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][31]  ( .D(n4523), .CP(n7256), .Q(
        \RegFilePlugin_regFile[9][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][31]  ( .D(n4491), .CP(n7191), .Q(
        \RegFilePlugin_regFile[8][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][31]  ( .D(n4459), .CP(n7239), .Q(
        \RegFilePlugin_regFile[7][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][31]  ( .D(n4427), .CP(n7256), .Q(
        \RegFilePlugin_regFile[6][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][31]  ( .D(n4395), .CP(n7256), .Q(
        \RegFilePlugin_regFile[5][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][31]  ( .D(n4363), .CP(n7239), .Q(
        \RegFilePlugin_regFile[4][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][31]  ( .D(n4331), .CP(n7239), .Q(
        \RegFilePlugin_regFile[3][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][31]  ( .D(n4299), .CP(n7192), .Q(
        \RegFilePlugin_regFile[2][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][31]  ( .D(n4267), .CP(n7239), .Q(
        \RegFilePlugin_regFile[1][31] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][31]  ( .D(n4234), .CP(n7192), .Q(
        \RegFilePlugin_regFile[0][31] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[31]  ( .D(N823), .CP(n7238), .Q(
        _zz_RegFilePlugin_regFile_port0[31]) );
  dfnrq1 \decode_to_execute_RS1_reg[31]  ( .D(n4233), .CP(n7193), .Q(
        execute_RS1[31]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[31]  ( .D(N856), .CP(n7239), .Q(
        _zz_RegFilePlugin_regFile_port1[31]) );
  dfnrq1 \decode_to_execute_RS2_reg[31]  ( .D(n4232), .CP(n7239), .Q(
        execute_RS2[31]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[31]  ( .D(
        n6206), .CP(n7238), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[31]) );
  dfnrq1 \CsrPlugin_mtval_reg[31]  ( .D(n6038), .CP(n7195), .Q(
        CsrPlugin_mtval[31]) );
  dfnrq1 \CsrPlugin_mepc_reg[31]  ( .D(n4080), .CP(n7188), .Q(
        CsrPlugin_mepc[31]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[31]  ( .D(n6164), .CP(
        n7239), .Q(_zz_CsrPlugin_csrMapping_readDataInit[31]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[30]  ( .D(N857), .CP(n7238), .Q(
        _zz_RegFilePlugin_regFile_port1[30]) );
  dfnrq1 \decode_to_execute_RS2_reg[30]  ( .D(n4229), .CP(n7239), .Q(
        execute_RS2[30]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][29]  ( .D(n5225), .CP(n7187), .Q(
        \RegFilePlugin_regFile[31][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][29]  ( .D(n5193), .CP(n7239), .Q(
        \RegFilePlugin_regFile[30][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][29]  ( .D(n5161), .CP(n7239), .Q(
        \RegFilePlugin_regFile[29][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][29]  ( .D(n5129), .CP(n7189), .Q(
        \RegFilePlugin_regFile[28][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][29]  ( .D(n5097), .CP(n7191), .Q(
        \RegFilePlugin_regFile[27][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][29]  ( .D(n5065), .CP(n7194), .Q(
        \RegFilePlugin_regFile[26][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][29]  ( .D(n5033), .CP(n7195), .Q(
        \RegFilePlugin_regFile[25][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][29]  ( .D(n5001), .CP(n7189), .Q(
        \RegFilePlugin_regFile[24][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][29]  ( .D(n4969), .CP(n7191), .Q(
        \RegFilePlugin_regFile[23][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][29]  ( .D(n4937), .CP(n7193), .Q(
        \RegFilePlugin_regFile[22][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][29]  ( .D(n4905), .CP(n7193), .Q(
        \RegFilePlugin_regFile[21][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][29]  ( .D(n4873), .CP(n7193), .Q(
        \RegFilePlugin_regFile[20][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][29]  ( .D(n4841), .CP(n7193), .Q(
        \RegFilePlugin_regFile[19][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][29]  ( .D(n4809), .CP(n7193), .Q(
        \RegFilePlugin_regFile[18][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][29]  ( .D(n4777), .CP(n7193), .Q(
        \RegFilePlugin_regFile[17][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][29]  ( .D(n4745), .CP(n7193), .Q(
        \RegFilePlugin_regFile[16][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][29]  ( .D(n4713), .CP(n7193), .Q(
        \RegFilePlugin_regFile[15][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][29]  ( .D(n4681), .CP(n7192), .Q(
        \RegFilePlugin_regFile[14][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][29]  ( .D(n4649), .CP(n7192), .Q(
        \RegFilePlugin_regFile[13][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][29]  ( .D(n4617), .CP(n7192), .Q(
        \RegFilePlugin_regFile[12][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][29]  ( .D(n4585), .CP(n7192), .Q(
        \RegFilePlugin_regFile[11][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][29]  ( .D(n4553), .CP(n7192), .Q(
        \RegFilePlugin_regFile[10][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][29]  ( .D(n4521), .CP(n7192), .Q(
        \RegFilePlugin_regFile[9][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][29]  ( .D(n4489), .CP(n7192), .Q(
        \RegFilePlugin_regFile[8][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][29]  ( .D(n4457), .CP(n7192), .Q(
        \RegFilePlugin_regFile[7][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][29]  ( .D(n4425), .CP(n7191), .Q(
        \RegFilePlugin_regFile[6][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][29]  ( .D(n4393), .CP(n7191), .Q(
        \RegFilePlugin_regFile[5][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][29]  ( .D(n4361), .CP(n7191), .Q(
        \RegFilePlugin_regFile[4][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][29]  ( .D(n4329), .CP(n7191), .Q(
        \RegFilePlugin_regFile[3][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][29]  ( .D(n4297), .CP(n7191), .Q(
        \RegFilePlugin_regFile[2][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][29]  ( .D(n4265), .CP(n7191), .Q(
        \RegFilePlugin_regFile[1][29] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][29]  ( .D(n4228), .CP(n7191), .Q(
        \RegFilePlugin_regFile[0][29] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[29]  ( .D(N825), .CP(n7191), .Q(
        _zz_RegFilePlugin_regFile_port0[29]) );
  dfnrq1 \decode_to_execute_RS1_reg[29]  ( .D(n4227), .CP(n7195), .Q(
        execute_RS1[29]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[29]  ( .D(n6162), .CP(
        n7188), .Q(_zz_CsrPlugin_csrMapping_readDataInit[29]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[27]  ( .D(n4114), .CP(n7192), .Q(
        CsrPlugin_mtvec_base[27]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[29]  ( .D(n6090), .CP(n7256), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[29]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[29]  ( .D(n5913), .CP(
        n7238), .Q(iBusWishbone_ADR[27]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[29]  ( 
        .D(n5312), .CP(n7194), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[29]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[29]  ( .D(
        n6204), .CP(n7193), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[29]) );
  dfnrq1 \CsrPlugin_mtval_reg[29]  ( .D(n6036), .CP(n7187), .Q(
        CsrPlugin_mtval[29]) );
  dfnrq1 \decode_to_execute_PC_reg[29]  ( .D(n5311), .CP(n7190), .Q(
        execute_PC[29]) );
  dfnrq1 \memory_to_writeBack_PC_reg[29]  ( .D(n5310), .CP(n7190), .Q(
        writeBack_PC[29]) );
  dfnrq1 \CsrPlugin_mepc_reg[29]  ( .D(n4082), .CP(n7190), .Q(
        CsrPlugin_mepc[29]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[29]  ( .D(n6043), .CP(n7190), .Q(
        debug_bus_rsp_data[29]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[29]  ( .D(N858), .CP(n7190), .Q(
        _zz_RegFilePlugin_regFile_port1[29]) );
  dfnrq1 \decode_to_execute_RS2_reg[29]  ( .D(n4226), .CP(n7190), .Q(
        execute_RS2[29]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][28]  ( .D(n5224), .CP(n7190), .Q(
        \RegFilePlugin_regFile[31][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][28]  ( .D(n5192), .CP(n7190), .Q(
        \RegFilePlugin_regFile[30][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][28]  ( .D(n5160), .CP(n7238), .Q(
        \RegFilePlugin_regFile[29][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][28]  ( .D(n5128), .CP(n7192), .Q(
        \RegFilePlugin_regFile[28][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][28]  ( .D(n5096), .CP(n7188), .Q(
        \RegFilePlugin_regFile[27][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][28]  ( .D(n5064), .CP(n7188), .Q(
        \RegFilePlugin_regFile[26][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][28]  ( .D(n5032), .CP(n7187), .Q(
        \RegFilePlugin_regFile[25][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][28]  ( .D(n5000), .CP(n7194), .Q(
        \RegFilePlugin_regFile[24][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][28]  ( .D(n4968), .CP(n7193), .Q(
        \RegFilePlugin_regFile[23][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][28]  ( .D(n4936), .CP(n7189), .Q(
        \RegFilePlugin_regFile[22][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][28]  ( .D(n4904), .CP(n7195), .Q(
        \RegFilePlugin_regFile[21][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][28]  ( .D(n4872), .CP(n7192), .Q(
        \RegFilePlugin_regFile[20][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][28]  ( .D(n4840), .CP(n7256), .Q(
        \RegFilePlugin_regFile[19][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][28]  ( .D(n4808), .CP(n7188), .Q(
        \RegFilePlugin_regFile[18][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][28]  ( .D(n4776), .CP(n7187), .Q(
        \RegFilePlugin_regFile[17][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][28]  ( .D(n4744), .CP(n7194), .Q(
        \RegFilePlugin_regFile[16][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][28]  ( .D(n4712), .CP(n7193), .Q(
        \RegFilePlugin_regFile[15][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][28]  ( .D(n4680), .CP(n7189), .Q(
        \RegFilePlugin_regFile[14][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][28]  ( .D(n4648), .CP(n7190), .Q(
        \RegFilePlugin_regFile[13][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][28]  ( .D(n4616), .CP(n7193), .Q(
        \RegFilePlugin_regFile[12][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][28]  ( .D(n4584), .CP(n7194), .Q(
        \RegFilePlugin_regFile[11][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][28]  ( .D(n4552), .CP(n7187), .Q(
        \RegFilePlugin_regFile[10][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][28]  ( .D(n4520), .CP(n7188), .Q(
        \RegFilePlugin_regFile[9][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][28]  ( .D(n4488), .CP(n7192), .Q(
        \RegFilePlugin_regFile[8][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][28]  ( .D(n4456), .CP(n7239), .Q(
        \RegFilePlugin_regFile[7][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][28]  ( .D(n4424), .CP(n7193), .Q(
        \RegFilePlugin_regFile[6][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][28]  ( .D(n4392), .CP(n7189), .Q(
        \RegFilePlugin_regFile[5][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][28]  ( .D(n4360), .CP(n7189), .Q(
        \RegFilePlugin_regFile[4][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][28]  ( .D(n4328), .CP(n7189), .Q(
        \RegFilePlugin_regFile[3][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][28]  ( .D(n4296), .CP(n7189), .Q(
        \RegFilePlugin_regFile[2][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][28]  ( .D(n4264), .CP(n7189), .Q(
        \RegFilePlugin_regFile[1][28] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][28]  ( .D(n4225), .CP(n7189), .Q(
        \RegFilePlugin_regFile[0][28] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[28]  ( .D(N826), .CP(n7189), .Q(
        _zz_RegFilePlugin_regFile_port0[28]) );
  dfnrq1 \decode_to_execute_RS1_reg[28]  ( .D(n4224), .CP(n7189), .Q(
        execute_RS1[28]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[28]  ( .D(n6161), .CP(
        n7188), .Q(_zz_CsrPlugin_csrMapping_readDataInit[28]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[26]  ( .D(n4115), .CP(n7188), .Q(
        CsrPlugin_mtvec_base[26]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[28]  ( .D(n6091), .CP(n7188), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[28]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[28]  ( .D(n5912), .CP(
        n7188), .Q(iBusWishbone_ADR[26]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[28]  ( 
        .D(n5309), .CP(n7188), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[28]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[28]  ( .D(
        n6203), .CP(n7188), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[28]) );
  dfnrq1 \CsrPlugin_mtval_reg[28]  ( .D(n6035), .CP(n7188), .Q(
        CsrPlugin_mtval[28]) );
  dfnrq1 \decode_to_execute_PC_reg[28]  ( .D(n5308), .CP(n7188), .Q(
        execute_PC[28]) );
  dfnrq1 \memory_to_writeBack_PC_reg[28]  ( .D(n5307), .CP(n7187), .Q(
        writeBack_PC[28]) );
  dfnrq1 \CsrPlugin_mepc_reg[28]  ( .D(n4083), .CP(n7190), .Q(
        CsrPlugin_mepc[28]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[28]  ( .D(n6044), .CP(n7194), .Q(
        debug_bus_rsp_data[28]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[28]  ( .D(N859), .CP(n7190), .Q(
        _zz_RegFilePlugin_regFile_port1[28]) );
  dfnrq1 \decode_to_execute_RS2_reg[28]  ( .D(n4223), .CP(n7193), .Q(
        execute_RS2[28]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][27]  ( .D(n5223), .CP(n7190), .Q(
        \RegFilePlugin_regFile[31][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][27]  ( .D(n5191), .CP(n7189), .Q(
        \RegFilePlugin_regFile[30][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][27]  ( .D(n5159), .CP(n7190), .Q(
        \RegFilePlugin_regFile[29][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][27]  ( .D(n5127), .CP(n7187), .Q(
        \RegFilePlugin_regFile[28][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][27]  ( .D(n5095), .CP(n7187), .Q(
        \RegFilePlugin_regFile[27][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][27]  ( .D(n5063), .CP(n7187), .Q(
        \RegFilePlugin_regFile[26][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][27]  ( .D(n5031), .CP(n7187), .Q(
        \RegFilePlugin_regFile[25][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][27]  ( .D(n4999), .CP(n7187), .Q(
        \RegFilePlugin_regFile[24][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][27]  ( .D(n4967), .CP(n7187), .Q(
        \RegFilePlugin_regFile[23][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][27]  ( .D(n4935), .CP(n7187), .Q(
        \RegFilePlugin_regFile[22][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][27]  ( .D(n4903), .CP(n7187), .Q(
        \RegFilePlugin_regFile[21][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][27]  ( .D(n4871), .CP(n7178), .Q(
        \RegFilePlugin_regFile[20][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][27]  ( .D(n4839), .CP(n7185), .Q(
        \RegFilePlugin_regFile[19][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][27]  ( .D(n4807), .CP(n7184), .Q(
        \RegFilePlugin_regFile[18][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][27]  ( .D(n4775), .CP(n7180), .Q(
        \RegFilePlugin_regFile[17][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][27]  ( .D(n4743), .CP(n7182), .Q(
        \RegFilePlugin_regFile[16][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][27]  ( .D(n4711), .CP(n7241), .Q(
        \RegFilePlugin_regFile[15][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][27]  ( .D(n4679), .CP(n7186), .Q(
        \RegFilePlugin_regFile[14][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][27]  ( .D(n4647), .CP(n7240), .Q(
        \RegFilePlugin_regFile[13][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][27]  ( .D(n4615), .CP(n7184), .Q(
        \RegFilePlugin_regFile[12][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][27]  ( .D(n4583), .CP(n7185), .Q(
        \RegFilePlugin_regFile[11][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][27]  ( .D(n4551), .CP(n7257), .Q(
        \RegFilePlugin_regFile[10][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][27]  ( .D(n4519), .CP(n7240), .Q(
        \RegFilePlugin_regFile[9][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][27]  ( .D(n4487), .CP(n7183), .Q(
        \RegFilePlugin_regFile[8][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][27]  ( .D(n4455), .CP(n7183), .Q(
        \RegFilePlugin_regFile[7][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][27]  ( .D(n4423), .CP(n7179), .Q(
        \RegFilePlugin_regFile[6][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][27]  ( .D(n4391), .CP(n7178), .Q(
        \RegFilePlugin_regFile[5][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][27]  ( .D(n4359), .CP(n7257), .Q(
        \RegFilePlugin_regFile[4][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][27]  ( .D(n4327), .CP(n7185), .Q(
        \RegFilePlugin_regFile[3][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][27]  ( .D(n4295), .CP(n7184), .Q(
        \RegFilePlugin_regFile[2][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][27]  ( .D(n4263), .CP(n7257), .Q(
        \RegFilePlugin_regFile[1][27] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][27]  ( .D(n4222), .CP(n7185), .Q(
        \RegFilePlugin_regFile[0][27] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[27]  ( .D(N827), .CP(n7257), .Q(
        _zz_RegFilePlugin_regFile_port0[27]) );
  dfnrq1 \decode_to_execute_RS1_reg[27]  ( .D(n4221), .CP(n7240), .Q(
        execute_RS1[27]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[27]  ( .D(n6160), .CP(
        n7183), .Q(_zz_CsrPlugin_csrMapping_readDataInit[27]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[25]  ( .D(n4116), .CP(n7183), .Q(
        CsrPlugin_mtvec_base[25]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[27]  ( .D(n6092), .CP(n7179), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[27]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[27]  ( .D(n5911), .CP(
        n7240), .Q(iBusWishbone_ADR[25]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[27]  ( 
        .D(n5306), .CP(n7182), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[27]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[27]  ( .D(
        n6202), .CP(n7178), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[27]) );
  dfnrq1 \CsrPlugin_mtval_reg[27]  ( .D(n6034), .CP(n7257), .Q(
        CsrPlugin_mtval[27]) );
  dfnrq1 \decode_to_execute_PC_reg[27]  ( .D(n5305), .CP(n7179), .Q(
        execute_PC[27]) );
  dfnrq1 \memory_to_writeBack_PC_reg[27]  ( .D(n5304), .CP(n7181), .Q(
        writeBack_PC[27]) );
  dfnrq1 \CsrPlugin_mepc_reg[27]  ( .D(n4084), .CP(n7240), .Q(
        CsrPlugin_mepc[27]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[27]  ( .D(n6045), .CP(n7240), .Q(
        debug_bus_rsp_data[27]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[27]  ( .D(N860), .CP(n7240), .Q(
        _zz_RegFilePlugin_regFile_port1[27]) );
  dfnrq1 \decode_to_execute_RS2_reg[27]  ( .D(n4220), .CP(n7240), .Q(
        execute_RS2[27]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][26]  ( .D(n5222), .CP(n7181), .Q(
        \RegFilePlugin_regFile[31][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][26]  ( .D(n5190), .CP(n7185), .Q(
        \RegFilePlugin_regFile[30][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][26]  ( .D(n5158), .CP(n7240), .Q(
        \RegFilePlugin_regFile[29][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][26]  ( .D(n5126), .CP(n7178), .Q(
        \RegFilePlugin_regFile[28][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][26]  ( .D(n5094), .CP(n7240), .Q(
        \RegFilePlugin_regFile[27][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][26]  ( .D(n5062), .CP(n7240), .Q(
        \RegFilePlugin_regFile[26][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][26]  ( .D(n5030), .CP(n7181), .Q(
        \RegFilePlugin_regFile[25][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][26]  ( .D(n4998), .CP(n7179), .Q(
        \RegFilePlugin_regFile[24][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][26]  ( .D(n4966), .CP(n7240), .Q(
        \RegFilePlugin_regFile[23][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][26]  ( .D(n4934), .CP(n7181), .Q(
        \RegFilePlugin_regFile[22][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][26]  ( .D(n4902), .CP(n7179), .Q(
        \RegFilePlugin_regFile[21][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][26]  ( .D(n4870), .CP(n7178), .Q(
        \RegFilePlugin_regFile[20][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][26]  ( .D(n4838), .CP(n7186), .Q(
        \RegFilePlugin_regFile[19][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][26]  ( .D(n4806), .CP(n7186), .Q(
        \RegFilePlugin_regFile[18][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][26]  ( .D(n4774), .CP(n7186), .Q(
        \RegFilePlugin_regFile[17][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][26]  ( .D(n4742), .CP(n7186), .Q(
        \RegFilePlugin_regFile[16][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][26]  ( .D(n4710), .CP(n7186), .Q(
        \RegFilePlugin_regFile[15][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][26]  ( .D(n4678), .CP(n7186), .Q(
        \RegFilePlugin_regFile[14][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][26]  ( .D(n4646), .CP(n7186), .Q(
        \RegFilePlugin_regFile[13][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][26]  ( .D(n4614), .CP(n7186), .Q(
        \RegFilePlugin_regFile[12][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][26]  ( .D(n4582), .CP(n7185), .Q(
        \RegFilePlugin_regFile[11][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][26]  ( .D(n4550), .CP(n7185), .Q(
        \RegFilePlugin_regFile[10][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][26]  ( .D(n4518), .CP(n7185), .Q(
        \RegFilePlugin_regFile[9][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][26]  ( .D(n4486), .CP(n7185), .Q(
        \RegFilePlugin_regFile[8][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][26]  ( .D(n4454), .CP(n7185), .Q(
        \RegFilePlugin_regFile[7][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][26]  ( .D(n4422), .CP(n7185), .Q(
        \RegFilePlugin_regFile[6][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][26]  ( .D(n4390), .CP(n7185), .Q(
        \RegFilePlugin_regFile[5][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][26]  ( .D(n4358), .CP(n7185), .Q(
        \RegFilePlugin_regFile[4][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][26]  ( .D(n4326), .CP(n7182), .Q(
        \RegFilePlugin_regFile[3][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][26]  ( .D(n4294), .CP(n7182), .Q(
        \RegFilePlugin_regFile[2][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][26]  ( .D(n4262), .CP(n7182), .Q(
        \RegFilePlugin_regFile[1][26] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][26]  ( .D(n4219), .CP(n7241), .Q(
        \RegFilePlugin_regFile[0][26] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[26]  ( .D(N828), .CP(n7182), .Q(
        _zz_RegFilePlugin_regFile_port0[26]) );
  dfnrq1 \decode_to_execute_RS1_reg[26]  ( .D(n4218), .CP(n7241), .Q(
        execute_RS1[26]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[26]  ( .D(n6159), .CP(
        n7182), .Q(_zz_CsrPlugin_csrMapping_readDataInit[26]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[24]  ( .D(n4117), .CP(n7241), .Q(
        CsrPlugin_mtvec_base[24]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[26]  ( .D(n6093), .CP(n7180), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[26]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[26]  ( .D(n5910), .CP(
        n7180), .Q(iBusWishbone_ADR[24]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[26]  ( 
        .D(n5303), .CP(n7180), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[26]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[26]  ( .D(
        n6201), .CP(n7186), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[26]) );
  dfnrq1 \CsrPlugin_mtval_reg[26]  ( .D(n6033), .CP(n7180), .Q(
        CsrPlugin_mtval[26]) );
  dfnrq1 \decode_to_execute_PC_reg[26]  ( .D(n5302), .CP(n7186), .Q(
        execute_PC[26]) );
  dfnrq1 \memory_to_writeBack_PC_reg[26]  ( .D(n5301), .CP(n7180), .Q(
        writeBack_PC[26]) );
  dfnrq1 \CsrPlugin_mepc_reg[26]  ( .D(n4085), .CP(n7186), .Q(
        CsrPlugin_mepc[26]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[26]  ( .D(n6046), .CP(n7257), .Q(
        debug_bus_rsp_data[26]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[26]  ( .D(N861), .CP(n7184), .Q(
        _zz_RegFilePlugin_regFile_port1[26]) );
  dfnrq1 \decode_to_execute_RS2_reg[26]  ( .D(n4217), .CP(n7257), .Q(
        execute_RS2[26]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][25]  ( .D(n5221), .CP(n7241), .Q(
        \RegFilePlugin_regFile[31][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][25]  ( .D(n5189), .CP(n7257), .Q(
        \RegFilePlugin_regFile[30][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][25]  ( .D(n5157), .CP(n7257), .Q(
        \RegFilePlugin_regFile[29][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][25]  ( .D(n5125), .CP(n7257), .Q(
        \RegFilePlugin_regFile[28][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][25]  ( .D(n5093), .CP(n7186), .Q(
        \RegFilePlugin_regFile[27][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][25]  ( .D(n5061), .CP(n7257), .Q(
        \RegFilePlugin_regFile[26][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][25]  ( .D(n5029), .CP(n7257), .Q(
        \RegFilePlugin_regFile[25][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][25]  ( .D(n4997), .CP(n7257), .Q(
        \RegFilePlugin_regFile[24][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][25]  ( .D(n4965), .CP(n7257), .Q(
        \RegFilePlugin_regFile[23][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][25]  ( .D(n4933), .CP(n7182), .Q(
        \RegFilePlugin_regFile[22][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][25]  ( .D(n4901), .CP(n7241), .Q(
        \RegFilePlugin_regFile[21][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][25]  ( .D(n4869), .CP(n7257), .Q(
        \RegFilePlugin_regFile[20][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][25]  ( .D(n4837), .CP(n7257), .Q(
        \RegFilePlugin_regFile[19][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][25]  ( .D(n4805), .CP(n7241), .Q(
        \RegFilePlugin_regFile[18][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][25]  ( .D(n4773), .CP(n7241), .Q(
        \RegFilePlugin_regFile[17][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][25]  ( .D(n4741), .CP(n7183), .Q(
        \RegFilePlugin_regFile[16][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][25]  ( .D(n4709), .CP(n7241), .Q(
        \RegFilePlugin_regFile[15][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][25]  ( .D(n4677), .CP(n7183), .Q(
        \RegFilePlugin_regFile[14][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][25]  ( .D(n4645), .CP(n7240), .Q(
        \RegFilePlugin_regFile[13][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][25]  ( .D(n4613), .CP(n7184), .Q(
        \RegFilePlugin_regFile[12][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][25]  ( .D(n4581), .CP(n7241), .Q(
        \RegFilePlugin_regFile[11][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][25]  ( .D(n4549), .CP(n7241), .Q(
        \RegFilePlugin_regFile[10][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][25]  ( .D(n4517), .CP(n7240), .Q(
        \RegFilePlugin_regFile[9][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][25]  ( .D(n4485), .CP(n7186), .Q(
        \RegFilePlugin_regFile[8][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][25]  ( .D(n4453), .CP(n7179), .Q(
        \RegFilePlugin_regFile[7][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][25]  ( .D(n4421), .CP(n7241), .Q(
        \RegFilePlugin_regFile[6][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][25]  ( .D(n4389), .CP(n7240), .Q(
        \RegFilePlugin_regFile[5][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][25]  ( .D(n4357), .CP(n7241), .Q(
        \RegFilePlugin_regFile[4][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][25]  ( .D(n4325), .CP(n7178), .Q(
        \RegFilePlugin_regFile[3][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][25]  ( .D(n4293), .CP(n7241), .Q(
        \RegFilePlugin_regFile[2][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][25]  ( .D(n4261), .CP(n7241), .Q(
        \RegFilePlugin_regFile[1][25] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][25]  ( .D(n4216), .CP(n7180), .Q(
        \RegFilePlugin_regFile[0][25] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[25]  ( .D(N829), .CP(n7182), .Q(
        _zz_RegFilePlugin_regFile_port0[25]) );
  dfnrq1 \decode_to_execute_RS1_reg[25]  ( .D(n4215), .CP(n7185), .Q(
        execute_RS1[25]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[25]  ( .D(n6158), .CP(
        n7186), .Q(_zz_CsrPlugin_csrMapping_readDataInit[25]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[23]  ( .D(n4118), .CP(n7180), .Q(
        CsrPlugin_mtvec_base[23]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[25]  ( .D(n6094), .CP(n7182), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[25]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[25]  ( .D(n5909), .CP(
        n7184), .Q(iBusWishbone_ADR[23]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[25]  ( 
        .D(n5300), .CP(n7184), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[25]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[25]  ( .D(
        n6200), .CP(n7184), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[25]) );
  dfnrq1 \CsrPlugin_mtval_reg[25]  ( .D(n6032), .CP(n7184), .Q(
        CsrPlugin_mtval[25]) );
  dfnrq1 \decode_to_execute_PC_reg[25]  ( .D(n5299), .CP(n7184), .Q(
        execute_PC[25]) );
  dfnrq1 \memory_to_writeBack_PC_reg[25]  ( .D(n5298), .CP(n7184), .Q(
        writeBack_PC[25]) );
  dfnrq1 \CsrPlugin_mepc_reg[25]  ( .D(n4086), .CP(n7184), .Q(
        CsrPlugin_mepc[25]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[25]  ( .D(n6047), .CP(n7184), .Q(
        debug_bus_rsp_data[25]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[25]  ( .D(N862), .CP(n7183), .Q(
        _zz_RegFilePlugin_regFile_port1[25]) );
  dfnrq1 \decode_to_execute_RS2_reg[25]  ( .D(n4214), .CP(n7183), .Q(
        execute_RS2[25]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][24]  ( .D(n5220), .CP(n7183), .Q(
        \RegFilePlugin_regFile[31][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][24]  ( .D(n5188), .CP(n7183), .Q(
        \RegFilePlugin_regFile[30][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][24]  ( .D(n5156), .CP(n7183), .Q(
        \RegFilePlugin_regFile[29][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][24]  ( .D(n5124), .CP(n7183), .Q(
        \RegFilePlugin_regFile[28][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][24]  ( .D(n5092), .CP(n7183), .Q(
        \RegFilePlugin_regFile[27][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][24]  ( .D(n5060), .CP(n7183), .Q(
        \RegFilePlugin_regFile[26][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][24]  ( .D(n5028), .CP(n7182), .Q(
        \RegFilePlugin_regFile[25][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][24]  ( .D(n4996), .CP(n7182), .Q(
        \RegFilePlugin_regFile[24][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][24]  ( .D(n4964), .CP(n7182), .Q(
        \RegFilePlugin_regFile[23][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][24]  ( .D(n4932), .CP(n7182), .Q(
        \RegFilePlugin_regFile[22][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][24]  ( .D(n4900), .CP(n7182), .Q(
        \RegFilePlugin_regFile[21][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][24]  ( .D(n4868), .CP(n7182), .Q(
        \RegFilePlugin_regFile[20][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][24]  ( .D(n4836), .CP(n7182), .Q(
        \RegFilePlugin_regFile[19][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][24]  ( .D(n4804), .CP(n7182), .Q(
        \RegFilePlugin_regFile[18][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][24]  ( .D(n4772), .CP(n7186), .Q(
        \RegFilePlugin_regFile[17][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][24]  ( .D(n4740), .CP(n7179), .Q(
        \RegFilePlugin_regFile[16][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][24]  ( .D(n4708), .CP(n7183), .Q(
        \RegFilePlugin_regFile[15][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][24]  ( .D(n4676), .CP(n7257), .Q(
        \RegFilePlugin_regFile[14][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][24]  ( .D(n4644), .CP(n7240), .Q(
        \RegFilePlugin_regFile[13][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][24]  ( .D(n4612), .CP(n7185), .Q(
        \RegFilePlugin_regFile[12][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][24]  ( .D(n4580), .CP(n7184), .Q(
        \RegFilePlugin_regFile[11][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][24]  ( .D(n4548), .CP(n7178), .Q(
        \RegFilePlugin_regFile[10][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][24]  ( .D(n4516), .CP(n7181), .Q(
        \RegFilePlugin_regFile[9][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][24]  ( .D(n4484), .CP(n7181), .Q(
        \RegFilePlugin_regFile[8][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][24]  ( .D(n4452), .CP(n7181), .Q(
        \RegFilePlugin_regFile[7][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][24]  ( .D(n4420), .CP(n7181), .Q(
        \RegFilePlugin_regFile[6][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][24]  ( .D(n4388), .CP(n7181), .Q(
        \RegFilePlugin_regFile[5][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][24]  ( .D(n4356), .CP(n7181), .Q(
        \RegFilePlugin_regFile[4][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][24]  ( .D(n4324), .CP(n7181), .Q(
        \RegFilePlugin_regFile[3][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][24]  ( .D(n4292), .CP(n7181), .Q(
        \RegFilePlugin_regFile[2][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][24]  ( .D(n4260), .CP(n7240), .Q(
        \RegFilePlugin_regFile[1][24] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][24]  ( .D(n4213), .CP(n7183), .Q(
        \RegFilePlugin_regFile[0][24] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[24]  ( .D(N830), .CP(n7179), .Q(
        _zz_RegFilePlugin_regFile_port0[24]) );
  dfnrq1 \decode_to_execute_RS1_reg[24]  ( .D(n4212), .CP(n7179), .Q(
        execute_RS1[24]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[24]  ( .D(n6157), .CP(
        n7178), .Q(_zz_CsrPlugin_csrMapping_readDataInit[24]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[22]  ( .D(n4119), .CP(n7185), .Q(
        CsrPlugin_mtvec_base[22]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[24]  ( .D(n6095), .CP(n7184), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[24]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[24]  ( .D(n5908), .CP(
        n7180), .Q(iBusWishbone_ADR[22]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[24]  ( 
        .D(n5297), .CP(n7186), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[24]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[24]  ( .D(
        n6199), .CP(n7183), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[24]) );
  dfnrq1 \CsrPlugin_mtval_reg[24]  ( .D(n6031), .CP(n7257), .Q(
        CsrPlugin_mtval[24]) );
  dfnrq1 \decode_to_execute_PC_reg[24]  ( .D(n5296), .CP(n7179), .Q(
        execute_PC[24]) );
  dfnrq1 \memory_to_writeBack_PC_reg[24]  ( .D(n5295), .CP(n7178), .Q(
        writeBack_PC[24]) );
  dfnrq1 \CsrPlugin_mepc_reg[24]  ( .D(n4087), .CP(n7185), .Q(
        CsrPlugin_mepc[24]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[24]  ( .D(n6048), .CP(n7184), .Q(
        debug_bus_rsp_data[24]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[24]  ( .D(N863), .CP(n7180), .Q(
        _zz_RegFilePlugin_regFile_port1[24]) );
  dfnrq1 \decode_to_execute_RS2_reg[24]  ( .D(n4211), .CP(n7181), .Q(
        execute_RS2[24]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][23]  ( .D(n5219), .CP(n7184), .Q(
        \RegFilePlugin_regFile[31][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][23]  ( .D(n5187), .CP(n7185), .Q(
        \RegFilePlugin_regFile[30][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][23]  ( .D(n5155), .CP(n7178), .Q(
        \RegFilePlugin_regFile[29][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][23]  ( .D(n5123), .CP(n7179), .Q(
        \RegFilePlugin_regFile[28][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][23]  ( .D(n5091), .CP(n7183), .Q(
        \RegFilePlugin_regFile[27][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][23]  ( .D(n5059), .CP(n7241), .Q(
        \RegFilePlugin_regFile[26][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][23]  ( .D(n5027), .CP(n7184), .Q(
        \RegFilePlugin_regFile[25][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][23]  ( .D(n4995), .CP(n7180), .Q(
        \RegFilePlugin_regFile[24][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][23]  ( .D(n4963), .CP(n7180), .Q(
        \RegFilePlugin_regFile[23][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][23]  ( .D(n4931), .CP(n7180), .Q(
        \RegFilePlugin_regFile[22][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][23]  ( .D(n4899), .CP(n7180), .Q(
        \RegFilePlugin_regFile[21][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][23]  ( .D(n4867), .CP(n7180), .Q(
        \RegFilePlugin_regFile[20][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][23]  ( .D(n4835), .CP(n7180), .Q(
        \RegFilePlugin_regFile[19][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][23]  ( .D(n4803), .CP(n7180), .Q(
        \RegFilePlugin_regFile[18][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][23]  ( .D(n4771), .CP(n7180), .Q(
        \RegFilePlugin_regFile[17][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][23]  ( .D(n4739), .CP(n7179), .Q(
        \RegFilePlugin_regFile[16][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][23]  ( .D(n4707), .CP(n7179), .Q(
        \RegFilePlugin_regFile[15][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][23]  ( .D(n4675), .CP(n7179), .Q(
        \RegFilePlugin_regFile[14][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][23]  ( .D(n4643), .CP(n7179), .Q(
        \RegFilePlugin_regFile[13][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][23]  ( .D(n4611), .CP(n7179), .Q(
        \RegFilePlugin_regFile[12][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][23]  ( .D(n4579), .CP(n7179), .Q(
        \RegFilePlugin_regFile[11][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][23]  ( .D(n4547), .CP(n7179), .Q(
        \RegFilePlugin_regFile[10][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][23]  ( .D(n4515), .CP(n7179), .Q(
        \RegFilePlugin_regFile[9][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][23]  ( .D(n4483), .CP(n7178), .Q(
        \RegFilePlugin_regFile[8][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][23]  ( .D(n4451), .CP(n7181), .Q(
        \RegFilePlugin_regFile[7][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][23]  ( .D(n4419), .CP(n7185), .Q(
        \RegFilePlugin_regFile[6][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][23]  ( .D(n4387), .CP(n7181), .Q(
        \RegFilePlugin_regFile[5][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][23]  ( .D(n4355), .CP(n7184), .Q(
        \RegFilePlugin_regFile[4][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][23]  ( .D(n4323), .CP(n7181), .Q(
        \RegFilePlugin_regFile[3][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][23]  ( .D(n4291), .CP(n7180), .Q(
        \RegFilePlugin_regFile[2][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][23]  ( .D(n4259), .CP(n7181), .Q(
        \RegFilePlugin_regFile[1][23] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][23]  ( .D(n4210), .CP(n7178), .Q(
        \RegFilePlugin_regFile[0][23] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[23]  ( .D(N831), .CP(n7178), .Q(
        _zz_RegFilePlugin_regFile_port0[23]) );
  dfnrq1 \decode_to_execute_RS1_reg[23]  ( .D(n4209), .CP(n7178), .Q(
        execute_RS1[23]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[23]  ( .D(n6156), .CP(
        n7178), .Q(_zz_CsrPlugin_csrMapping_readDataInit[23]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[21]  ( .D(n4120), .CP(n7178), .Q(
        CsrPlugin_mtvec_base[21]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[23]  ( .D(n6096), .CP(n7178), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[23]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[23]  ( .D(n5907), .CP(
        n7178), .Q(iBusWishbone_ADR[21]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[23]  ( 
        .D(n5294), .CP(n7178), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[23]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[23]  ( .D(
        n6198), .CP(n7169), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[23]) );
  dfnrq1 \CsrPlugin_mtval_reg[23]  ( .D(n6030), .CP(n7176), .Q(
        CsrPlugin_mtval[23]) );
  dfnrq1 \decode_to_execute_PC_reg[23]  ( .D(n5293), .CP(n7175), .Q(
        execute_PC[23]) );
  dfnrq1 \memory_to_writeBack_PC_reg[23]  ( .D(n5292), .CP(n7171), .Q(
        writeBack_PC[23]) );
  dfnrq1 \CsrPlugin_mepc_reg[23]  ( .D(n4088), .CP(n7173), .Q(
        CsrPlugin_mepc[23]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[23]  ( .D(n6049), .CP(n7243), .Q(
        debug_bus_rsp_data[23]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[23]  ( .D(N864), .CP(n7177), .Q(
        _zz_RegFilePlugin_regFile_port1[23]) );
  dfnrq1 \decode_to_execute_RS2_reg[23]  ( .D(n4208), .CP(n7242), .Q(
        execute_RS2[23]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][22]  ( .D(n5218), .CP(n7175), .Q(
        \RegFilePlugin_regFile[31][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][22]  ( .D(n5186), .CP(n7176), .Q(
        \RegFilePlugin_regFile[30][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][22]  ( .D(n5154), .CP(n7258), .Q(
        \RegFilePlugin_regFile[29][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][22]  ( .D(n5122), .CP(n7242), .Q(
        \RegFilePlugin_regFile[28][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][22]  ( .D(n5090), .CP(n7174), .Q(
        \RegFilePlugin_regFile[27][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][22]  ( .D(n5058), .CP(n7174), .Q(
        \RegFilePlugin_regFile[26][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][22]  ( .D(n5026), .CP(n7170), .Q(
        \RegFilePlugin_regFile[25][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][22]  ( .D(n4994), .CP(n7169), .Q(
        \RegFilePlugin_regFile[24][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][22]  ( .D(n4962), .CP(n7258), .Q(
        \RegFilePlugin_regFile[23][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][22]  ( .D(n4930), .CP(n7176), .Q(
        \RegFilePlugin_regFile[22][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][22]  ( .D(n4898), .CP(n7175), .Q(
        \RegFilePlugin_regFile[21][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][22]  ( .D(n4866), .CP(n7258), .Q(
        \RegFilePlugin_regFile[20][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][22]  ( .D(n4834), .CP(n7176), .Q(
        \RegFilePlugin_regFile[19][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][22]  ( .D(n4802), .CP(n7258), .Q(
        \RegFilePlugin_regFile[18][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][22]  ( .D(n4770), .CP(n7242), .Q(
        \RegFilePlugin_regFile[17][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][22]  ( .D(n4738), .CP(n7174), .Q(
        \RegFilePlugin_regFile[16][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][22]  ( .D(n4706), .CP(n7174), .Q(
        \RegFilePlugin_regFile[15][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][22]  ( .D(n4674), .CP(n7170), .Q(
        \RegFilePlugin_regFile[14][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][22]  ( .D(n4642), .CP(n7242), .Q(
        \RegFilePlugin_regFile[13][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][22]  ( .D(n4610), .CP(n7173), .Q(
        \RegFilePlugin_regFile[12][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][22]  ( .D(n4578), .CP(n7169), .Q(
        \RegFilePlugin_regFile[11][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][22]  ( .D(n4546), .CP(n7258), .Q(
        \RegFilePlugin_regFile[10][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][22]  ( .D(n4514), .CP(n7170), .Q(
        \RegFilePlugin_regFile[9][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][22]  ( .D(n4482), .CP(n7172), .Q(
        \RegFilePlugin_regFile[8][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][22]  ( .D(n4450), .CP(n7242), .Q(
        \RegFilePlugin_regFile[7][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][22]  ( .D(n4418), .CP(n7242), .Q(
        \RegFilePlugin_regFile[6][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][22]  ( .D(n4386), .CP(n7242), .Q(
        \RegFilePlugin_regFile[5][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][22]  ( .D(n4354), .CP(n7242), .Q(
        \RegFilePlugin_regFile[4][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][22]  ( .D(n4322), .CP(n7172), .Q(
        \RegFilePlugin_regFile[3][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][22]  ( .D(n4290), .CP(n7176), .Q(
        \RegFilePlugin_regFile[2][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][22]  ( .D(n4258), .CP(n7242), .Q(
        \RegFilePlugin_regFile[1][22] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][22]  ( .D(n4207), .CP(n7169), .Q(
        \RegFilePlugin_regFile[0][22] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[22]  ( .D(N832), .CP(n7242), .Q(
        _zz_RegFilePlugin_regFile_port0[22]) );
  dfnrq1 \decode_to_execute_RS1_reg[22]  ( .D(n4206), .CP(n7242), .Q(
        execute_RS1[22]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[22]  ( .D(n6155), .CP(
        n7172), .Q(_zz_CsrPlugin_csrMapping_readDataInit[22]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[20]  ( .D(n4121), .CP(n7170), .Q(
        CsrPlugin_mtvec_base[20]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[22]  ( .D(n6097), .CP(n7242), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[22]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[22]  ( .D(n5906), .CP(
        n7172), .Q(iBusWishbone_ADR[20]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[22]  ( 
        .D(n5291), .CP(n7170), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[22]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[22]  ( .D(
        n6197), .CP(n7169), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[22]) );
  dfnrq1 \CsrPlugin_mtval_reg[22]  ( .D(n6029), .CP(n7177), .Q(
        CsrPlugin_mtval[22]) );
  dfnrq1 \decode_to_execute_PC_reg[22]  ( .D(n5290), .CP(n7177), .Q(
        execute_PC[22]) );
  dfnrq1 \memory_to_writeBack_PC_reg[22]  ( .D(n5289), .CP(n7177), .Q(
        writeBack_PC[22]) );
  dfnrq1 \CsrPlugin_mepc_reg[22]  ( .D(n4089), .CP(n7177), .Q(
        CsrPlugin_mepc[22]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[22]  ( .D(n6050), .CP(n7177), .Q(
        debug_bus_rsp_data[22]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[22]  ( .D(N865), .CP(n7177), .Q(
        _zz_RegFilePlugin_regFile_port1[22]) );
  dfnrq1 \decode_to_execute_RS2_reg[22]  ( .D(n4205), .CP(n7177), .Q(
        execute_RS2[22]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][21]  ( .D(n5217), .CP(n7177), .Q(
        \RegFilePlugin_regFile[31][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][21]  ( .D(n5185), .CP(n7176), .Q(
        \RegFilePlugin_regFile[30][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][21]  ( .D(n5153), .CP(n7176), .Q(
        \RegFilePlugin_regFile[29][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][21]  ( .D(n5121), .CP(n7176), .Q(
        \RegFilePlugin_regFile[28][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][21]  ( .D(n5089), .CP(n7176), .Q(
        \RegFilePlugin_regFile[27][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][21]  ( .D(n5057), .CP(n7176), .Q(
        \RegFilePlugin_regFile[26][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][21]  ( .D(n5025), .CP(n7176), .Q(
        \RegFilePlugin_regFile[25][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][21]  ( .D(n4993), .CP(n7176), .Q(
        \RegFilePlugin_regFile[24][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][21]  ( .D(n4961), .CP(n7176), .Q(
        \RegFilePlugin_regFile[23][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][21]  ( .D(n4929), .CP(n7173), .Q(
        \RegFilePlugin_regFile[22][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][21]  ( .D(n4897), .CP(n7173), .Q(
        \RegFilePlugin_regFile[21][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][21]  ( .D(n4865), .CP(n7173), .Q(
        \RegFilePlugin_regFile[20][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][21]  ( .D(n4833), .CP(n7243), .Q(
        \RegFilePlugin_regFile[19][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][21]  ( .D(n4801), .CP(n7173), .Q(
        \RegFilePlugin_regFile[18][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][21]  ( .D(n4769), .CP(n7243), .Q(
        \RegFilePlugin_regFile[17][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][21]  ( .D(n4737), .CP(n7173), .Q(
        \RegFilePlugin_regFile[16][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][21]  ( .D(n4705), .CP(n7243), .Q(
        \RegFilePlugin_regFile[15][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][21]  ( .D(n4673), .CP(n7171), .Q(
        \RegFilePlugin_regFile[14][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][21]  ( .D(n4641), .CP(n7171), .Q(
        \RegFilePlugin_regFile[13][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][21]  ( .D(n4609), .CP(n7171), .Q(
        \RegFilePlugin_regFile[12][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][21]  ( .D(n4577), .CP(n7177), .Q(
        \RegFilePlugin_regFile[11][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][21]  ( .D(n4545), .CP(n7171), .Q(
        \RegFilePlugin_regFile[10][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][21]  ( .D(n4513), .CP(n7177), .Q(
        \RegFilePlugin_regFile[9][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][21]  ( .D(n4481), .CP(n7171), .Q(
        \RegFilePlugin_regFile[8][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][21]  ( .D(n4449), .CP(n7177), .Q(
        \RegFilePlugin_regFile[7][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][21]  ( .D(n4417), .CP(n7258), .Q(
        \RegFilePlugin_regFile[6][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][21]  ( .D(n4385), .CP(n7175), .Q(
        \RegFilePlugin_regFile[5][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][21]  ( .D(n4353), .CP(n7258), .Q(
        \RegFilePlugin_regFile[4][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][21]  ( .D(n4321), .CP(n7243), .Q(
        \RegFilePlugin_regFile[3][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][21]  ( .D(n4289), .CP(n7258), .Q(
        \RegFilePlugin_regFile[2][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][21]  ( .D(n4257), .CP(n7258), .Q(
        \RegFilePlugin_regFile[1][21] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][21]  ( .D(n4204), .CP(n7258), .Q(
        \RegFilePlugin_regFile[0][21] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[21]  ( .D(N833), .CP(n7177), .Q(
        _zz_RegFilePlugin_regFile_port0[21]) );
  dfnrq1 \decode_to_execute_RS1_reg[21]  ( .D(n4203), .CP(n7258), .Q(
        execute_RS1[21]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[21]  ( .D(n6154), .CP(
        n7258), .Q(_zz_CsrPlugin_csrMapping_readDataInit[21]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[19]  ( .D(n4122), .CP(n7258), .Q(
        CsrPlugin_mtvec_base[19]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[21]  ( .D(n6098), .CP(n7258), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[21]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[21]  ( .D(n5905), .CP(
        n7173), .Q(iBusWishbone_ADR[19]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[21]  ( 
        .D(n5288), .CP(n7243), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[21]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[21]  ( .D(
        n6196), .CP(n7258), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[21]) );
  dfnrq1 \CsrPlugin_mtval_reg[21]  ( .D(n6028), .CP(n7258), .Q(
        CsrPlugin_mtval[21]) );
  dfnrq1 \decode_to_execute_PC_reg[21]  ( .D(n5287), .CP(n7243), .Q(
        execute_PC[21]) );
  dfnrq1 \memory_to_writeBack_PC_reg[21]  ( .D(n5286), .CP(n7243), .Q(
        writeBack_PC[21]) );
  dfnrq1 \CsrPlugin_mepc_reg[21]  ( .D(n4090), .CP(n7174), .Q(
        CsrPlugin_mepc[21]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[21]  ( .D(n6051), .CP(n7243), .Q(
        debug_bus_rsp_data[21]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[21]  ( .D(N866), .CP(n7174), .Q(
        _zz_RegFilePlugin_regFile_port1[21]) );
  dfnrq1 \decode_to_execute_RS2_reg[21]  ( .D(n4202), .CP(n7242), .Q(
        execute_RS2[21]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][20]  ( .D(n5216), .CP(n7175), .Q(
        \RegFilePlugin_regFile[31][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][20]  ( .D(n5184), .CP(n7243), .Q(
        \RegFilePlugin_regFile[30][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][20]  ( .D(n5152), .CP(n7243), .Q(
        \RegFilePlugin_regFile[29][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][20]  ( .D(n5120), .CP(n7242), .Q(
        \RegFilePlugin_regFile[28][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][20]  ( .D(n5088), .CP(n7177), .Q(
        \RegFilePlugin_regFile[27][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][20]  ( .D(n5056), .CP(n7170), .Q(
        \RegFilePlugin_regFile[26][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][20]  ( .D(n5024), .CP(n7243), .Q(
        \RegFilePlugin_regFile[25][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][20]  ( .D(n4992), .CP(n7242), .Q(
        \RegFilePlugin_regFile[24][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][20]  ( .D(n4960), .CP(n7243), .Q(
        \RegFilePlugin_regFile[23][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][20]  ( .D(n4928), .CP(n7169), .Q(
        \RegFilePlugin_regFile[22][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][20]  ( .D(n4896), .CP(n7243), .Q(
        \RegFilePlugin_regFile[21][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][20]  ( .D(n4864), .CP(n7243), .Q(
        \RegFilePlugin_regFile[20][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][20]  ( .D(n4832), .CP(n7171), .Q(
        \RegFilePlugin_regFile[19][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][20]  ( .D(n4800), .CP(n7173), .Q(
        \RegFilePlugin_regFile[18][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][20]  ( .D(n4768), .CP(n7176), .Q(
        \RegFilePlugin_regFile[17][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][20]  ( .D(n4736), .CP(n7177), .Q(
        \RegFilePlugin_regFile[16][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][20]  ( .D(n4704), .CP(n7171), .Q(
        \RegFilePlugin_regFile[15][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][20]  ( .D(n4672), .CP(n7173), .Q(
        \RegFilePlugin_regFile[14][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][20]  ( .D(n4640), .CP(n7175), .Q(
        \RegFilePlugin_regFile[13][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][20]  ( .D(n4608), .CP(n7175), .Q(
        \RegFilePlugin_regFile[12][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][20]  ( .D(n4576), .CP(n7175), .Q(
        \RegFilePlugin_regFile[11][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][20]  ( .D(n4544), .CP(n7175), .Q(
        \RegFilePlugin_regFile[10][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][20]  ( .D(n4512), .CP(n7175), .Q(
        \RegFilePlugin_regFile[9][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][20]  ( .D(n4480), .CP(n7175), .Q(
        \RegFilePlugin_regFile[8][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][20]  ( .D(n4448), .CP(n7175), .Q(
        \RegFilePlugin_regFile[7][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][20]  ( .D(n4416), .CP(n7175), .Q(
        \RegFilePlugin_regFile[6][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][20]  ( .D(n4384), .CP(n7174), .Q(
        \RegFilePlugin_regFile[5][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][20]  ( .D(n4352), .CP(n7174), .Q(
        \RegFilePlugin_regFile[4][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][20]  ( .D(n4320), .CP(n7174), .Q(
        \RegFilePlugin_regFile[3][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][20]  ( .D(n4288), .CP(n7174), .Q(
        \RegFilePlugin_regFile[2][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][20]  ( .D(n4256), .CP(n7174), .Q(
        \RegFilePlugin_regFile[1][20] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][20]  ( .D(n4201), .CP(n7174), .Q(
        \RegFilePlugin_regFile[0][20] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[20]  ( .D(N834), .CP(n7174), .Q(
        _zz_RegFilePlugin_regFile_port0[20]) );
  dfnrq1 \decode_to_execute_RS1_reg[20]  ( .D(n4200), .CP(n7174), .Q(
        execute_RS1[20]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[20]  ( .D(n6153), .CP(
        n7173), .Q(_zz_CsrPlugin_csrMapping_readDataInit[20]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[18]  ( .D(n4123), .CP(n7173), .Q(
        CsrPlugin_mtvec_base[18]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[20]  ( .D(n6099), .CP(n7173), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[20]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[20]  ( .D(n5904), .CP(
        n7173), .Q(iBusWishbone_ADR[18]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[20]  ( 
        .D(n5285), .CP(n7173), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[20]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[20]  ( .D(
        n6195), .CP(n7173), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[20]) );
  dfnrq1 \CsrPlugin_mtval_reg[20]  ( .D(n6027), .CP(n7173), .Q(
        CsrPlugin_mtval[20]) );
  dfnrq1 \decode_to_execute_PC_reg[20]  ( .D(n5284), .CP(n7173), .Q(
        execute_PC[20]) );
  dfnrq1 \memory_to_writeBack_PC_reg[20]  ( .D(n5283), .CP(n7177), .Q(
        writeBack_PC[20]) );
  dfnrq1 \CsrPlugin_mepc_reg[20]  ( .D(n4091), .CP(n7170), .Q(
        CsrPlugin_mepc[20]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[20]  ( .D(n6052), .CP(n7174), .Q(
        debug_bus_rsp_data[20]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[20]  ( .D(N867), .CP(n7258), .Q(
        _zz_RegFilePlugin_regFile_port1[20]) );
  dfnrq1 \decode_to_execute_RS2_reg[20]  ( .D(n4199), .CP(n7242), .Q(
        execute_RS2[20]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][19]  ( .D(n5215), .CP(n7176), .Q(
        \RegFilePlugin_regFile[31][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][19]  ( .D(n5183), .CP(n7175), .Q(
        \RegFilePlugin_regFile[30][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][19]  ( .D(n5151), .CP(n7169), .Q(
        \RegFilePlugin_regFile[29][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][19]  ( .D(n5119), .CP(n7172), .Q(
        \RegFilePlugin_regFile[28][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][19]  ( .D(n5087), .CP(n7172), .Q(
        \RegFilePlugin_regFile[27][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][19]  ( .D(n5055), .CP(n7172), .Q(
        \RegFilePlugin_regFile[26][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][19]  ( .D(n5023), .CP(n7172), .Q(
        \RegFilePlugin_regFile[25][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][19]  ( .D(n4991), .CP(n7172), .Q(
        \RegFilePlugin_regFile[24][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][19]  ( .D(n4959), .CP(n7172), .Q(
        \RegFilePlugin_regFile[23][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][19]  ( .D(n4927), .CP(n7172), .Q(
        \RegFilePlugin_regFile[22][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][19]  ( .D(n4895), .CP(n7172), .Q(
        \RegFilePlugin_regFile[21][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][19]  ( .D(n4863), .CP(n7242), .Q(
        \RegFilePlugin_regFile[20][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][19]  ( .D(n4831), .CP(n7174), .Q(
        \RegFilePlugin_regFile[19][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][19]  ( .D(n4799), .CP(n7170), .Q(
        \RegFilePlugin_regFile[18][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][19]  ( .D(n4767), .CP(n7170), .Q(
        \RegFilePlugin_regFile[17][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][19]  ( .D(n4735), .CP(n7169), .Q(
        \RegFilePlugin_regFile[16][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][19]  ( .D(n4703), .CP(n7176), .Q(
        \RegFilePlugin_regFile[15][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][19]  ( .D(n4671), .CP(n7175), .Q(
        \RegFilePlugin_regFile[14][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][19]  ( .D(n4639), .CP(n7171), .Q(
        \RegFilePlugin_regFile[13][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][19]  ( .D(n4607), .CP(n7177), .Q(
        \RegFilePlugin_regFile[12][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][19]  ( .D(n4575), .CP(n7174), .Q(
        \RegFilePlugin_regFile[11][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][19]  ( .D(n4543), .CP(n7258), .Q(
        \RegFilePlugin_regFile[10][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][19]  ( .D(n4511), .CP(n7170), .Q(
        \RegFilePlugin_regFile[9][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][19]  ( .D(n4479), .CP(n7169), .Q(
        \RegFilePlugin_regFile[8][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][19]  ( .D(n4447), .CP(n7176), .Q(
        \RegFilePlugin_regFile[7][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][19]  ( .D(n4415), .CP(n7175), .Q(
        \RegFilePlugin_regFile[6][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][19]  ( .D(n4383), .CP(n7171), .Q(
        \RegFilePlugin_regFile[5][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][19]  ( .D(n4351), .CP(n7172), .Q(
        \RegFilePlugin_regFile[4][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][19]  ( .D(n4319), .CP(n7175), .Q(
        \RegFilePlugin_regFile[3][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][19]  ( .D(n4287), .CP(n7176), .Q(
        \RegFilePlugin_regFile[2][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][19]  ( .D(n4255), .CP(n7169), .Q(
        \RegFilePlugin_regFile[1][19] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][19]  ( .D(n4198), .CP(n7170), .Q(
        \RegFilePlugin_regFile[0][19] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[19]  ( .D(N835), .CP(n7174), .Q(
        _zz_RegFilePlugin_regFile_port0[19]) );
  dfnrq1 \decode_to_execute_RS1_reg[19]  ( .D(n4197), .CP(n7243), .Q(
        execute_RS1[19]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[19]  ( .D(n6152), .CP(
        n7175), .Q(_zz_CsrPlugin_csrMapping_readDataInit[19]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[17]  ( .D(n4124), .CP(n7171), .Q(
        CsrPlugin_mtvec_base[17]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[19]  ( .D(n6100), .CP(n7171), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[19]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[19]  ( .D(n5903), .CP(
        n7171), .Q(iBusWishbone_ADR[17]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[19]  ( 
        .D(n5282), .CP(n7171), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[19]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[19]  ( .D(
        n6194), .CP(n7171), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[19]) );
  dfnrq1 \CsrPlugin_mtval_reg[19]  ( .D(n6026), .CP(n7171), .Q(
        CsrPlugin_mtval[19]) );
  dfnrq1 \decode_to_execute_PC_reg[19]  ( .D(n5281), .CP(n7171), .Q(
        execute_PC[19]) );
  dfnrq1 \memory_to_writeBack_PC_reg[19]  ( .D(n5280), .CP(n7171), .Q(
        writeBack_PC[19]) );
  dfnrq1 \CsrPlugin_mepc_reg[19]  ( .D(n4092), .CP(n7170), .Q(
        CsrPlugin_mepc[19]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[19]  ( .D(n6053), .CP(n7170), .Q(
        debug_bus_rsp_data[19]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[19]  ( .D(N868), .CP(n7170), .Q(
        _zz_RegFilePlugin_regFile_port1[19]) );
  dfnrq1 \decode_to_execute_RS2_reg[19]  ( .D(n4196), .CP(n7170), .Q(
        execute_RS2[19]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][18]  ( .D(n5214), .CP(n7170), .Q(
        \RegFilePlugin_regFile[31][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][18]  ( .D(n5182), .CP(n7170), .Q(
        \RegFilePlugin_regFile[30][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][18]  ( .D(n5150), .CP(n7170), .Q(
        \RegFilePlugin_regFile[29][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][18]  ( .D(n5118), .CP(n7170), .Q(
        \RegFilePlugin_regFile[28][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][18]  ( .D(n5086), .CP(n7169), .Q(
        \RegFilePlugin_regFile[27][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][18]  ( .D(n5054), .CP(n7172), .Q(
        \RegFilePlugin_regFile[26][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][18]  ( .D(n5022), .CP(n7176), .Q(
        \RegFilePlugin_regFile[25][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][18]  ( .D(n4990), .CP(n7172), .Q(
        \RegFilePlugin_regFile[24][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][18]  ( .D(n4958), .CP(n7175), .Q(
        \RegFilePlugin_regFile[23][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][18]  ( .D(n4926), .CP(n7172), .Q(
        \RegFilePlugin_regFile[22][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][18]  ( .D(n4894), .CP(n7171), .Q(
        \RegFilePlugin_regFile[21][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][18]  ( .D(n4862), .CP(n7172), .Q(
        \RegFilePlugin_regFile[20][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][18]  ( .D(n4830), .CP(n7169), .Q(
        \RegFilePlugin_regFile[19][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][18]  ( .D(n4798), .CP(n7169), .Q(
        \RegFilePlugin_regFile[18][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][18]  ( .D(n4766), .CP(n7169), .Q(
        \RegFilePlugin_regFile[17][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][18]  ( .D(n4734), .CP(n7169), .Q(
        \RegFilePlugin_regFile[16][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][18]  ( .D(n4702), .CP(n7169), .Q(
        \RegFilePlugin_regFile[15][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][18]  ( .D(n4670), .CP(n7169), .Q(
        \RegFilePlugin_regFile[14][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][18]  ( .D(n4638), .CP(n7169), .Q(
        \RegFilePlugin_regFile[13][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][18]  ( .D(n4606), .CP(n7169), .Q(
        \RegFilePlugin_regFile[12][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][18]  ( .D(n4574), .CP(n7160), .Q(
        \RegFilePlugin_regFile[11][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][18]  ( .D(n4542), .CP(n7167), .Q(
        \RegFilePlugin_regFile[10][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][18]  ( .D(n4510), .CP(n7166), .Q(
        \RegFilePlugin_regFile[9][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][18]  ( .D(n4478), .CP(n7162), .Q(
        \RegFilePlugin_regFile[8][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][18]  ( .D(n4446), .CP(n7164), .Q(
        \RegFilePlugin_regFile[7][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][18]  ( .D(n4414), .CP(n7245), .Q(
        \RegFilePlugin_regFile[6][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][18]  ( .D(n4382), .CP(n7168), .Q(
        \RegFilePlugin_regFile[5][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][18]  ( .D(n4350), .CP(n7244), .Q(
        \RegFilePlugin_regFile[4][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][18]  ( .D(n4318), .CP(n7166), .Q(
        \RegFilePlugin_regFile[3][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][18]  ( .D(n4286), .CP(n7167), .Q(
        \RegFilePlugin_regFile[2][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][18]  ( .D(n4254), .CP(n7259), .Q(
        \RegFilePlugin_regFile[1][18] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][18]  ( .D(n4195), .CP(n7244), .Q(
        \RegFilePlugin_regFile[0][18] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[18]  ( .D(N836), .CP(n7165), .Q(
        _zz_RegFilePlugin_regFile_port0[18]) );
  dfnrq1 \decode_to_execute_RS1_reg[18]  ( .D(n4194), .CP(n7165), .Q(
        execute_RS1[18]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[18]  ( .D(n6151), .CP(
        n7161), .Q(_zz_CsrPlugin_csrMapping_readDataInit[18]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[16]  ( .D(n4125), .CP(n7160), .Q(
        CsrPlugin_mtvec_base[16]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[18]  ( .D(n6101), .CP(n7259), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[18]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[18]  ( .D(n5902), .CP(
        n7167), .Q(iBusWishbone_ADR[16]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[18]  ( 
        .D(n5279), .CP(n7166), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[18]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[18]  ( .D(
        n6193), .CP(n7259), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[18]) );
  dfnrq1 \CsrPlugin_mtval_reg[18]  ( .D(n6025), .CP(n7167), .Q(
        CsrPlugin_mtval[18]) );
  dfnrq1 \decode_to_execute_PC_reg[18]  ( .D(n5278), .CP(n7259), .Q(
        execute_PC[18]) );
  dfnrq1 \memory_to_writeBack_PC_reg[18]  ( .D(n5277), .CP(n7244), .Q(
        writeBack_PC[18]) );
  dfnrq1 \CsrPlugin_mepc_reg[18]  ( .D(n4093), .CP(n7165), .Q(
        CsrPlugin_mepc[18]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[18]  ( .D(n6054), .CP(n7165), .Q(
        debug_bus_rsp_data[18]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[18]  ( .D(N869), .CP(n7161), .Q(
        _zz_RegFilePlugin_regFile_port1[18]) );
  dfnrq1 \decode_to_execute_RS2_reg[18]  ( .D(n4193), .CP(n7244), .Q(
        execute_RS2[18]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][17]  ( .D(n5213), .CP(n7164), .Q(
        \RegFilePlugin_regFile[31][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][17]  ( .D(n5181), .CP(n7160), .Q(
        \RegFilePlugin_regFile[30][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][17]  ( .D(n5149), .CP(n7259), .Q(
        \RegFilePlugin_regFile[29][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][17]  ( .D(n5117), .CP(n7161), .Q(
        \RegFilePlugin_regFile[28][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][17]  ( .D(n5085), .CP(n7163), .Q(
        \RegFilePlugin_regFile[27][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][17]  ( .D(n5053), .CP(n7244), .Q(
        \RegFilePlugin_regFile[26][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][17]  ( .D(n5021), .CP(n7244), .Q(
        \RegFilePlugin_regFile[25][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][17]  ( .D(n4989), .CP(n7244), .Q(
        \RegFilePlugin_regFile[24][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][17]  ( .D(n4957), .CP(n7244), .Q(
        \RegFilePlugin_regFile[23][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][17]  ( .D(n4925), .CP(n7163), .Q(
        \RegFilePlugin_regFile[22][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][17]  ( .D(n4893), .CP(n7167), .Q(
        \RegFilePlugin_regFile[21][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][17]  ( .D(n4861), .CP(n7244), .Q(
        \RegFilePlugin_regFile[20][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][17]  ( .D(n4829), .CP(n7160), .Q(
        \RegFilePlugin_regFile[19][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][17]  ( .D(n4797), .CP(n7244), .Q(
        \RegFilePlugin_regFile[18][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][17]  ( .D(n4765), .CP(n7244), .Q(
        \RegFilePlugin_regFile[17][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][17]  ( .D(n4733), .CP(n7163), .Q(
        \RegFilePlugin_regFile[16][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][17]  ( .D(n4701), .CP(n7161), .Q(
        \RegFilePlugin_regFile[15][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][17]  ( .D(n4669), .CP(n7244), .Q(
        \RegFilePlugin_regFile[14][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][17]  ( .D(n4637), .CP(n7163), .Q(
        \RegFilePlugin_regFile[13][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][17]  ( .D(n4605), .CP(n7161), .Q(
        \RegFilePlugin_regFile[12][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][17]  ( .D(n4573), .CP(n7160), .Q(
        \RegFilePlugin_regFile[11][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][17]  ( .D(n4541), .CP(n7168), .Q(
        \RegFilePlugin_regFile[10][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][17]  ( .D(n4509), .CP(n7168), .Q(
        \RegFilePlugin_regFile[9][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][17]  ( .D(n4477), .CP(n7168), .Q(
        \RegFilePlugin_regFile[8][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][17]  ( .D(n4445), .CP(n7168), .Q(
        \RegFilePlugin_regFile[7][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][17]  ( .D(n4413), .CP(n7168), .Q(
        \RegFilePlugin_regFile[6][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][17]  ( .D(n4381), .CP(n7168), .Q(
        \RegFilePlugin_regFile[5][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][17]  ( .D(n4349), .CP(n7168), .Q(
        \RegFilePlugin_regFile[4][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][17]  ( .D(n4317), .CP(n7168), .Q(
        \RegFilePlugin_regFile[3][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][17]  ( .D(n4285), .CP(n7167), .Q(
        \RegFilePlugin_regFile[2][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][17]  ( .D(n4253), .CP(n7167), .Q(
        \RegFilePlugin_regFile[1][17] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][17]  ( .D(n4192), .CP(n7167), .Q(
        \RegFilePlugin_regFile[0][17] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[17]  ( .D(N837), .CP(n7167), .Q(
        _zz_RegFilePlugin_regFile_port0[17]) );
  dfnrq1 \decode_to_execute_RS1_reg[17]  ( .D(n4191), .CP(n7167), .Q(
        execute_RS1[17]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[17]  ( .D(n6150), .CP(
        n7167), .Q(_zz_CsrPlugin_csrMapping_readDataInit[17]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[15]  ( .D(n4126), .CP(n7167), .Q(
        CsrPlugin_mtvec_base[15]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[17]  ( .D(n6102), .CP(n7167), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[17]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[17]  ( .D(n5901), .CP(
        n7164), .Q(iBusWishbone_ADR[15]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[17]  ( 
        .D(n5276), .CP(n7164), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[17]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[17]  ( .D(
        n6192), .CP(n7164), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[17]) );
  dfnrq1 \CsrPlugin_mtval_reg[17]  ( .D(n6024), .CP(n7245), .Q(
        CsrPlugin_mtval[17]) );
  dfnrq1 \decode_to_execute_PC_reg[17]  ( .D(n5275), .CP(n7164), .Q(
        execute_PC[17]) );
  dfnrq1 \memory_to_writeBack_PC_reg[17]  ( .D(n5274), .CP(n7245), .Q(
        writeBack_PC[17]) );
  dfnrq1 \CsrPlugin_mepc_reg[17]  ( .D(n4094), .CP(n7164), .Q(
        CsrPlugin_mepc[17]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[17]  ( .D(n6055), .CP(n7245), .Q(
        debug_bus_rsp_data[17]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[17]  ( .D(N870), .CP(n7162), .Q(
        _zz_RegFilePlugin_regFile_port1[17]) );
  dfnrq1 \decode_to_execute_RS2_reg[17]  ( .D(n4190), .CP(n7162), .Q(
        execute_RS2[17]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][16]  ( .D(n5212), .CP(n7162), .Q(
        \RegFilePlugin_regFile[31][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][16]  ( .D(n5180), .CP(n7168), .Q(
        \RegFilePlugin_regFile[30][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][16]  ( .D(n5148), .CP(n7162), .Q(
        \RegFilePlugin_regFile[29][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][16]  ( .D(n5116), .CP(n7168), .Q(
        \RegFilePlugin_regFile[28][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][16]  ( .D(n5084), .CP(n7162), .Q(
        \RegFilePlugin_regFile[27][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][16]  ( .D(n5052), .CP(n7168), .Q(
        \RegFilePlugin_regFile[26][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][16]  ( .D(n5020), .CP(n7259), .Q(
        \RegFilePlugin_regFile[25][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][16]  ( .D(n4988), .CP(n7166), .Q(
        \RegFilePlugin_regFile[24][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][16]  ( .D(n4956), .CP(n7259), .Q(
        \RegFilePlugin_regFile[23][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][16]  ( .D(n4924), .CP(n7245), .Q(
        \RegFilePlugin_regFile[22][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][16]  ( .D(n4892), .CP(n7259), .Q(
        \RegFilePlugin_regFile[21][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][16]  ( .D(n4860), .CP(n7259), .Q(
        \RegFilePlugin_regFile[20][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][16]  ( .D(n4828), .CP(n7259), .Q(
        \RegFilePlugin_regFile[19][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][16]  ( .D(n4796), .CP(n7168), .Q(
        \RegFilePlugin_regFile[18][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][16]  ( .D(n4764), .CP(n7259), .Q(
        \RegFilePlugin_regFile[17][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][16]  ( .D(n4732), .CP(n7259), .Q(
        \RegFilePlugin_regFile[16][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][16]  ( .D(n4700), .CP(n7259), .Q(
        \RegFilePlugin_regFile[15][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][16]  ( .D(n4668), .CP(n7259), .Q(
        \RegFilePlugin_regFile[14][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][16]  ( .D(n4636), .CP(n7164), .Q(
        \RegFilePlugin_regFile[13][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][16]  ( .D(n4604), .CP(n7245), .Q(
        \RegFilePlugin_regFile[12][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][16]  ( .D(n4572), .CP(n7259), .Q(
        \RegFilePlugin_regFile[11][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][16]  ( .D(n4540), .CP(n7259), .Q(
        \RegFilePlugin_regFile[10][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][16]  ( .D(n4508), .CP(n7245), .Q(
        \RegFilePlugin_regFile[9][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][16]  ( .D(n4476), .CP(n7245), .Q(
        \RegFilePlugin_regFile[8][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][16]  ( .D(n4444), .CP(n7165), .Q(
        \RegFilePlugin_regFile[7][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][16]  ( .D(n4412), .CP(n7245), .Q(
        \RegFilePlugin_regFile[6][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][16]  ( .D(n4380), .CP(n7165), .Q(
        \RegFilePlugin_regFile[5][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][16]  ( .D(n4348), .CP(n7244), .Q(
        \RegFilePlugin_regFile[4][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][16]  ( .D(n4316), .CP(n7166), .Q(
        \RegFilePlugin_regFile[3][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][16]  ( .D(n4284), .CP(n7245), .Q(
        \RegFilePlugin_regFile[2][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][16]  ( .D(n4252), .CP(n7245), .Q(
        \RegFilePlugin_regFile[1][16] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][16]  ( .D(n4189), .CP(n7244), .Q(
        \RegFilePlugin_regFile[0][16] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[16]  ( .D(N838), .CP(n7168), .Q(
        _zz_RegFilePlugin_regFile_port0[16]) );
  dfnrq1 \decode_to_execute_RS1_reg[16]  ( .D(n4188), .CP(n7161), .Q(
        execute_RS1[16]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[16]  ( .D(n6149), .CP(
        n7245), .Q(_zz_CsrPlugin_csrMapping_readDataInit[16]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[14]  ( .D(n4127), .CP(n7244), .Q(
        CsrPlugin_mtvec_base[14]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[16]  ( .D(n6103), .CP(n7245), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[16]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[16]  ( .D(n5900), .CP(
        n7160), .Q(iBusWishbone_ADR[14]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[16]  ( 
        .D(n5273), .CP(n7245), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[16]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[16]  ( .D(
        n6191), .CP(n7245), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[16]) );
  dfnrq1 \CsrPlugin_mtval_reg[16]  ( .D(n6023), .CP(n7162), .Q(
        CsrPlugin_mtval[16]) );
  dfnrq1 \decode_to_execute_PC_reg[16]  ( .D(n5272), .CP(n7164), .Q(
        execute_PC[16]) );
  dfnrq1 \memory_to_writeBack_PC_reg[16]  ( .D(n5271), .CP(n7167), .Q(
        writeBack_PC[16]) );
  dfnrq1 \CsrPlugin_mepc_reg[16]  ( .D(n4095), .CP(n7168), .Q(
        CsrPlugin_mepc[16]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[16]  ( .D(n6056), .CP(n7162), .Q(
        debug_bus_rsp_data[16]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[16]  ( .D(N871), .CP(n7164), .Q(
        _zz_RegFilePlugin_regFile_port1[16]) );
  dfnrq1 \decode_to_execute_RS2_reg[16]  ( .D(n4187), .CP(n7166), .Q(
        execute_RS2[16]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][15]  ( .D(n5211), .CP(n7166), .Q(
        \RegFilePlugin_regFile[31][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][15]  ( .D(n5179), .CP(n7166), .Q(
        \RegFilePlugin_regFile[30][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][15]  ( .D(n5147), .CP(n7166), .Q(
        \RegFilePlugin_regFile[29][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][15]  ( .D(n5115), .CP(n7166), .Q(
        \RegFilePlugin_regFile[28][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][15]  ( .D(n5083), .CP(n7166), .Q(
        \RegFilePlugin_regFile[27][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][15]  ( .D(n5051), .CP(n7166), .Q(
        \RegFilePlugin_regFile[26][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][15]  ( .D(n5019), .CP(n7166), .Q(
        \RegFilePlugin_regFile[25][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][15]  ( .D(n4987), .CP(n7165), .Q(
        \RegFilePlugin_regFile[24][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][15]  ( .D(n4955), .CP(n7165), .Q(
        \RegFilePlugin_regFile[23][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][15]  ( .D(n4923), .CP(n7165), .Q(
        \RegFilePlugin_regFile[22][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][15]  ( .D(n4891), .CP(n7165), .Q(
        \RegFilePlugin_regFile[21][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][15]  ( .D(n4859), .CP(n7165), .Q(
        \RegFilePlugin_regFile[20][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][15]  ( .D(n4827), .CP(n7165), .Q(
        \RegFilePlugin_regFile[19][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][15]  ( .D(n4795), .CP(n7165), .Q(
        \RegFilePlugin_regFile[18][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][15]  ( .D(n4763), .CP(n7165), .Q(
        \RegFilePlugin_regFile[17][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][15]  ( .D(n4731), .CP(n7164), .Q(
        \RegFilePlugin_regFile[16][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][15]  ( .D(n4699), .CP(n7164), .Q(
        \RegFilePlugin_regFile[15][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][15]  ( .D(n4667), .CP(n7164), .Q(
        \RegFilePlugin_regFile[14][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][15]  ( .D(n4635), .CP(n7164), .Q(
        \RegFilePlugin_regFile[13][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][15]  ( .D(n4603), .CP(n7164), .Q(
        \RegFilePlugin_regFile[12][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][15]  ( .D(n4571), .CP(n7164), .Q(
        \RegFilePlugin_regFile[11][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][15]  ( .D(n4539), .CP(n7164), .Q(
        \RegFilePlugin_regFile[10][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][15]  ( .D(n4507), .CP(n7164), .Q(
        \RegFilePlugin_regFile[9][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][15]  ( .D(n4475), .CP(n7168), .Q(
        \RegFilePlugin_regFile[8][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][15]  ( .D(n4443), .CP(n7161), .Q(
        \RegFilePlugin_regFile[7][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][15]  ( .D(n4411), .CP(n7165), .Q(
        \RegFilePlugin_regFile[6][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][15]  ( .D(n4379), .CP(n7259), .Q(
        \RegFilePlugin_regFile[5][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][15]  ( .D(n4347), .CP(n7244), .Q(
        \RegFilePlugin_regFile[4][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][15]  ( .D(n4315), .CP(n7167), .Q(
        \RegFilePlugin_regFile[3][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][15]  ( .D(n4283), .CP(n7166), .Q(
        \RegFilePlugin_regFile[2][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][15]  ( .D(n4251), .CP(n7160), .Q(
        \RegFilePlugin_regFile[1][15] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][15]  ( .D(n4186), .CP(n7163), .Q(
        \RegFilePlugin_regFile[0][15] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[15]  ( .D(N839), .CP(n7163), .Q(
        _zz_RegFilePlugin_regFile_port0[15]) );
  dfnrq1 \decode_to_execute_RS1_reg[15]  ( .D(n4185), .CP(n7163), .Q(
        execute_RS1[15]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[15]  ( .D(n6148), .CP(
        n7163), .Q(_zz_CsrPlugin_csrMapping_readDataInit[15]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[13]  ( .D(n4128), .CP(n7163), .Q(
        CsrPlugin_mtvec_base[13]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[15]  ( .D(n6104), .CP(n7163), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[15]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[15]  ( .D(n5899), .CP(
        n7163), .Q(iBusWishbone_ADR[13]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[15]  ( 
        .D(n5270), .CP(n7163), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[15]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[15]  ( .D(
        n6190), .CP(n7244), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[15]) );
  dfnrq1 \CsrPlugin_mtval_reg[15]  ( .D(n6022), .CP(n7165), .Q(
        CsrPlugin_mtval[15]) );
  dfnrq1 \decode_to_execute_PC_reg[15]  ( .D(n5269), .CP(n7161), .Q(
        execute_PC[15]) );
  dfnrq1 \memory_to_writeBack_PC_reg[15]  ( .D(n5268), .CP(n7161), .Q(
        writeBack_PC[15]) );
  dfnrq1 \CsrPlugin_mepc_reg[15]  ( .D(n4096), .CP(n7160), .Q(
        CsrPlugin_mepc[15]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[15]  ( .D(n6057), .CP(n7167), .Q(
        debug_bus_rsp_data[15]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[15]  ( .D(N872), .CP(n7166), .Q(
        _zz_RegFilePlugin_regFile_port1[15]) );
  dfnrq1 \decode_to_execute_RS2_reg[15]  ( .D(n4184), .CP(n7162), .Q(
        execute_RS2[15]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][14]  ( .D(n5210), .CP(n7168), .Q(
        \RegFilePlugin_regFile[31][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][14]  ( .D(n5178), .CP(n7165), .Q(
        \RegFilePlugin_regFile[30][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][14]  ( .D(n5146), .CP(n7259), .Q(
        \RegFilePlugin_regFile[29][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][14]  ( .D(n5114), .CP(n7161), .Q(
        \RegFilePlugin_regFile[28][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][14]  ( .D(n5082), .CP(n7160), .Q(
        \RegFilePlugin_regFile[27][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][14]  ( .D(n5050), .CP(n7167), .Q(
        \RegFilePlugin_regFile[26][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][14]  ( .D(n5018), .CP(n7166), .Q(
        \RegFilePlugin_regFile[25][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][14]  ( .D(n4986), .CP(n7162), .Q(
        \RegFilePlugin_regFile[24][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][14]  ( .D(n4954), .CP(n7163), .Q(
        \RegFilePlugin_regFile[23][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][14]  ( .D(n4922), .CP(n7166), .Q(
        \RegFilePlugin_regFile[22][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][14]  ( .D(n4890), .CP(n7167), .Q(
        \RegFilePlugin_regFile[21][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][14]  ( .D(n4858), .CP(n7160), .Q(
        \RegFilePlugin_regFile[20][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][14]  ( .D(n4826), .CP(n7161), .Q(
        \RegFilePlugin_regFile[19][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][14]  ( .D(n4794), .CP(n7165), .Q(
        \RegFilePlugin_regFile[18][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][14]  ( .D(n4762), .CP(n7245), .Q(
        \RegFilePlugin_regFile[17][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][14]  ( .D(n4730), .CP(n7166), .Q(
        \RegFilePlugin_regFile[16][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][14]  ( .D(n4698), .CP(n7162), .Q(
        \RegFilePlugin_regFile[15][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][14]  ( .D(n4666), .CP(n7162), .Q(
        \RegFilePlugin_regFile[14][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][14]  ( .D(n4634), .CP(n7162), .Q(
        \RegFilePlugin_regFile[13][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][14]  ( .D(n4602), .CP(n7162), .Q(
        \RegFilePlugin_regFile[12][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][14]  ( .D(n4570), .CP(n7162), .Q(
        \RegFilePlugin_regFile[11][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][14]  ( .D(n4538), .CP(n7162), .Q(
        \RegFilePlugin_regFile[10][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][14]  ( .D(n4506), .CP(n7162), .Q(
        \RegFilePlugin_regFile[9][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][14]  ( .D(n4474), .CP(n7162), .Q(
        \RegFilePlugin_regFile[8][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][14]  ( .D(n4442), .CP(n7161), .Q(
        \RegFilePlugin_regFile[7][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][14]  ( .D(n4410), .CP(n7161), .Q(
        \RegFilePlugin_regFile[6][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][14]  ( .D(n4378), .CP(n7161), .Q(
        \RegFilePlugin_regFile[5][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][14]  ( .D(n4346), .CP(n7161), .Q(
        \RegFilePlugin_regFile[4][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][14]  ( .D(n4314), .CP(n7161), .Q(
        \RegFilePlugin_regFile[3][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][14]  ( .D(n4282), .CP(n7161), .Q(
        \RegFilePlugin_regFile[2][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][14]  ( .D(n4250), .CP(n7161), .Q(
        \RegFilePlugin_regFile[1][14] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][14]  ( .D(n4183), .CP(n7161), .Q(
        \RegFilePlugin_regFile[0][14] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[14]  ( .D(N840), .CP(n7160), .Q(
        _zz_RegFilePlugin_regFile_port0[14]) );
  dfnrq1 \decode_to_execute_RS1_reg[14]  ( .D(n4182), .CP(n7163), .Q(
        execute_RS1[14]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[14]  ( .D(n6147), .CP(
        n7167), .Q(_zz_CsrPlugin_csrMapping_readDataInit[14]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[12]  ( .D(n4129), .CP(n7163), .Q(
        CsrPlugin_mtvec_base[12]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[14]  ( .D(n6105), .CP(n7166), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[14]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[14]  ( .D(n5898), .CP(
        n7163), .Q(iBusWishbone_ADR[12]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[14]  ( 
        .D(n5267), .CP(n7162), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[14]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[14]  ( .D(
        n6189), .CP(n7163), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[14]) );
  dfnrq1 \CsrPlugin_mtval_reg[14]  ( .D(n6021), .CP(n7160), .Q(
        CsrPlugin_mtval[14]) );
  dfnrq1 \decode_to_execute_PC_reg[14]  ( .D(n5266), .CP(n7160), .Q(
        execute_PC[14]) );
  dfnrq1 \memory_to_writeBack_PC_reg[14]  ( .D(n5265), .CP(n7160), .Q(
        writeBack_PC[14]) );
  dfnrq1 \CsrPlugin_mepc_reg[14]  ( .D(n4097), .CP(n7160), .Q(
        CsrPlugin_mepc[14]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[14]  ( .D(n6058), .CP(n7160), .Q(
        debug_bus_rsp_data[14]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[14]  ( .D(N873), .CP(n7160), .Q(
        _zz_RegFilePlugin_regFile_port1[14]) );
  dfnrq1 \decode_to_execute_RS2_reg[14]  ( .D(n4181), .CP(n7160), .Q(
        execute_RS2[14]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][13]  ( .D(n5209), .CP(n7160), .Q(
        \RegFilePlugin_regFile[31][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][13]  ( .D(n5177), .CP(n7151), .Q(
        \RegFilePlugin_regFile[30][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][13]  ( .D(n5145), .CP(n7158), .Q(
        \RegFilePlugin_regFile[29][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][13]  ( .D(n5113), .CP(n7157), .Q(
        \RegFilePlugin_regFile[28][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][13]  ( .D(n5081), .CP(n7153), .Q(
        \RegFilePlugin_regFile[27][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][13]  ( .D(n5049), .CP(n7155), .Q(
        \RegFilePlugin_regFile[26][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][13]  ( .D(n5017), .CP(n7247), .Q(
        \RegFilePlugin_regFile[25][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][13]  ( .D(n4985), .CP(n7159), .Q(
        \RegFilePlugin_regFile[24][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][13]  ( .D(n4953), .CP(n7246), .Q(
        \RegFilePlugin_regFile[23][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][13]  ( .D(n4921), .CP(n7157), .Q(
        \RegFilePlugin_regFile[22][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][13]  ( .D(n4889), .CP(n7158), .Q(
        \RegFilePlugin_regFile[21][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][13]  ( .D(n4857), .CP(n7260), .Q(
        \RegFilePlugin_regFile[20][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][13]  ( .D(n4825), .CP(n7246), .Q(
        \RegFilePlugin_regFile[19][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][13]  ( .D(n4793), .CP(n7156), .Q(
        \RegFilePlugin_regFile[18][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][13]  ( .D(n4761), .CP(n7156), .Q(
        \RegFilePlugin_regFile[17][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][13]  ( .D(n4729), .CP(n7152), .Q(
        \RegFilePlugin_regFile[16][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][13]  ( .D(n4697), .CP(n7151), .Q(
        \RegFilePlugin_regFile[15][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][13]  ( .D(n4665), .CP(n7260), .Q(
        \RegFilePlugin_regFile[14][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][13]  ( .D(n4633), .CP(n7158), .Q(
        \RegFilePlugin_regFile[13][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][13]  ( .D(n4601), .CP(n7157), .Q(
        \RegFilePlugin_regFile[12][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][13]  ( .D(n4569), .CP(n7260), .Q(
        \RegFilePlugin_regFile[11][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][13]  ( .D(n4537), .CP(n7158), .Q(
        \RegFilePlugin_regFile[10][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][13]  ( .D(n4505), .CP(n7260), .Q(
        \RegFilePlugin_regFile[9][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][13]  ( .D(n4473), .CP(n7246), .Q(
        \RegFilePlugin_regFile[8][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][13]  ( .D(n4441), .CP(n7156), .Q(
        \RegFilePlugin_regFile[7][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][13]  ( .D(n4409), .CP(n7156), .Q(
        \RegFilePlugin_regFile[6][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][13]  ( .D(n4377), .CP(n7152), .Q(
        \RegFilePlugin_regFile[5][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][13]  ( .D(n4345), .CP(n7246), .Q(
        \RegFilePlugin_regFile[4][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][13]  ( .D(n4313), .CP(n7155), .Q(
        \RegFilePlugin_regFile[3][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][13]  ( .D(n4281), .CP(n7151), .Q(
        \RegFilePlugin_regFile[2][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][13]  ( .D(n4249), .CP(n7260), .Q(
        \RegFilePlugin_regFile[1][13] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][13]  ( .D(n4180), .CP(n7152), .Q(
        \RegFilePlugin_regFile[0][13] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[13]  ( .D(N841), .CP(n7154), .Q(
        _zz_RegFilePlugin_regFile_port0[13]) );
  dfnrq1 \decode_to_execute_RS1_reg[13]  ( .D(n4179), .CP(n7246), .Q(
        execute_RS1[13]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[13]  ( .D(n6146), .CP(
        n7246), .Q(_zz_CsrPlugin_csrMapping_readDataInit[13]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[11]  ( .D(n4130), .CP(n7246), .Q(
        CsrPlugin_mtvec_base[11]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[13]  ( .D(n6106), .CP(n7246), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[13]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[13]  ( .D(n5897), .CP(
        n7154), .Q(iBusWishbone_ADR[11]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[13]  ( 
        .D(n5264), .CP(n7158), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[13]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[13]  ( .D(
        n6188), .CP(n7246), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[13]) );
  dfnrq1 \CsrPlugin_mtval_reg[13]  ( .D(n6020), .CP(n7151), .Q(
        CsrPlugin_mtval[13]) );
  dfnrq1 \decode_to_execute_PC_reg[13]  ( .D(n5263), .CP(n7246), .Q(
        execute_PC[13]) );
  dfnrq1 \memory_to_writeBack_PC_reg[13]  ( .D(n5262), .CP(n7246), .Q(
        writeBack_PC[13]) );
  dfnrq1 \CsrPlugin_mepc_reg[13]  ( .D(n4098), .CP(n7154), .Q(
        CsrPlugin_mepc[13]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[13]  ( .D(n6059), .CP(n7152), .Q(
        debug_bus_rsp_data[13]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[13]  ( .D(N874), .CP(n7246), .Q(
        _zz_RegFilePlugin_regFile_port1[13]) );
  dfnrq1 \decode_to_execute_RS2_reg[13]  ( .D(n4178), .CP(n7154), .Q(
        execute_RS2[13]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][12]  ( .D(n5208), .CP(n7152), .Q(
        \RegFilePlugin_regFile[31][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][12]  ( .D(n5176), .CP(n7151), .Q(
        \RegFilePlugin_regFile[30][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][12]  ( .D(n5144), .CP(n7159), .Q(
        \RegFilePlugin_regFile[29][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][12]  ( .D(n5112), .CP(n7159), .Q(
        \RegFilePlugin_regFile[28][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][12]  ( .D(n5080), .CP(n7159), .Q(
        \RegFilePlugin_regFile[27][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][12]  ( .D(n5048), .CP(n7159), .Q(
        \RegFilePlugin_regFile[26][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][12]  ( .D(n5016), .CP(n7159), .Q(
        \RegFilePlugin_regFile[25][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][12]  ( .D(n4984), .CP(n7159), .Q(
        \RegFilePlugin_regFile[24][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][12]  ( .D(n4952), .CP(n7159), .Q(
        \RegFilePlugin_regFile[23][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][12]  ( .D(n4920), .CP(n7159), .Q(
        \RegFilePlugin_regFile[22][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][12]  ( .D(n4888), .CP(n7158), .Q(
        \RegFilePlugin_regFile[21][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][12]  ( .D(n4856), .CP(n7158), .Q(
        \RegFilePlugin_regFile[20][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][12]  ( .D(n4824), .CP(n7158), .Q(
        \RegFilePlugin_regFile[19][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][12]  ( .D(n4792), .CP(n7158), .Q(
        \RegFilePlugin_regFile[18][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][12]  ( .D(n4760), .CP(n7158), .Q(
        \RegFilePlugin_regFile[17][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][12]  ( .D(n4728), .CP(n7158), .Q(
        \RegFilePlugin_regFile[16][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][12]  ( .D(n4696), .CP(n7158), .Q(
        \RegFilePlugin_regFile[15][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][12]  ( .D(n4664), .CP(n7158), .Q(
        \RegFilePlugin_regFile[14][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][12]  ( .D(n4632), .CP(n7155), .Q(
        \RegFilePlugin_regFile[13][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][12]  ( .D(n4600), .CP(n7155), .Q(
        \RegFilePlugin_regFile[12][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][12]  ( .D(n4568), .CP(n7155), .Q(
        \RegFilePlugin_regFile[11][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][12]  ( .D(n4536), .CP(n7247), .Q(
        \RegFilePlugin_regFile[10][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][12]  ( .D(n4504), .CP(n7155), .Q(
        \RegFilePlugin_regFile[9][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][12]  ( .D(n4472), .CP(n7247), .Q(
        \RegFilePlugin_regFile[8][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][12]  ( .D(n4440), .CP(n7155), .Q(
        \RegFilePlugin_regFile[7][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][12]  ( .D(n4408), .CP(n7247), .Q(
        \RegFilePlugin_regFile[6][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][12]  ( .D(n4376), .CP(n7153), .Q(
        \RegFilePlugin_regFile[5][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][12]  ( .D(n4344), .CP(n7153), .Q(
        \RegFilePlugin_regFile[4][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][12]  ( .D(n4312), .CP(n7153), .Q(
        \RegFilePlugin_regFile[3][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][12]  ( .D(n4280), .CP(n7159), .Q(
        \RegFilePlugin_regFile[2][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][12]  ( .D(n4248), .CP(n7153), .Q(
        \RegFilePlugin_regFile[1][12] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][12]  ( .D(n4177), .CP(n7159), .Q(
        \RegFilePlugin_regFile[0][12] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[12]  ( .D(N842), .CP(n7153), .Q(
        _zz_RegFilePlugin_regFile_port0[12]) );
  dfnrq1 \decode_to_execute_RS1_reg[12]  ( .D(n4176), .CP(n7159), .Q(
        execute_RS1[12]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[12]  ( .D(N875), .CP(n7260), .Q(
        _zz_RegFilePlugin_regFile_port1[12]) );
  dfnrq1 \decode_to_execute_RS2_reg[12]  ( .D(n4175), .CP(n7157), .Q(
        execute_RS2[12]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][11]  ( .D(n5207), .CP(n7260), .Q(
        \RegFilePlugin_regFile[31][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][11]  ( .D(n5175), .CP(n7247), .Q(
        \RegFilePlugin_regFile[30][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][11]  ( .D(n5143), .CP(n7260), .Q(
        \RegFilePlugin_regFile[29][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][11]  ( .D(n5111), .CP(n7260), .Q(
        \RegFilePlugin_regFile[28][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][11]  ( .D(n5079), .CP(n7260), .Q(
        \RegFilePlugin_regFile[27][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][11]  ( .D(n5047), .CP(n7159), .Q(
        \RegFilePlugin_regFile[26][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][11]  ( .D(n5015), .CP(n7260), .Q(
        \RegFilePlugin_regFile[25][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][11]  ( .D(n4983), .CP(n7260), .Q(
        \RegFilePlugin_regFile[24][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][11]  ( .D(n4951), .CP(n7260), .Q(
        \RegFilePlugin_regFile[23][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][11]  ( .D(n4919), .CP(n7260), .Q(
        \RegFilePlugin_regFile[22][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][11]  ( .D(n4887), .CP(n7155), .Q(
        \RegFilePlugin_regFile[21][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][11]  ( .D(n4855), .CP(n7247), .Q(
        \RegFilePlugin_regFile[20][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][11]  ( .D(n4823), .CP(n7260), .Q(
        \RegFilePlugin_regFile[19][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][11]  ( .D(n4791), .CP(n7260), .Q(
        \RegFilePlugin_regFile[18][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][11]  ( .D(n4759), .CP(n7247), .Q(
        \RegFilePlugin_regFile[17][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][11]  ( .D(n4727), .CP(n7247), .Q(
        \RegFilePlugin_regFile[16][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][11]  ( .D(n4695), .CP(n7156), .Q(
        \RegFilePlugin_regFile[15][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][11]  ( .D(n4663), .CP(n7247), .Q(
        \RegFilePlugin_regFile[14][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][11]  ( .D(n4631), .CP(n7156), .Q(
        \RegFilePlugin_regFile[13][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][11]  ( .D(n4599), .CP(n7246), .Q(
        \RegFilePlugin_regFile[12][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][11]  ( .D(n4567), .CP(n7157), .Q(
        \RegFilePlugin_regFile[11][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][11]  ( .D(n4535), .CP(n7247), .Q(
        \RegFilePlugin_regFile[10][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][11]  ( .D(n4503), .CP(n7247), .Q(
        \RegFilePlugin_regFile[9][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][11]  ( .D(n4471), .CP(n7246), .Q(
        \RegFilePlugin_regFile[8][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][11]  ( .D(n4439), .CP(n7159), .Q(
        \RegFilePlugin_regFile[7][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][11]  ( .D(n4407), .CP(n7152), .Q(
        \RegFilePlugin_regFile[6][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][11]  ( .D(n4375), .CP(n7247), .Q(
        \RegFilePlugin_regFile[5][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][11]  ( .D(n4343), .CP(n7246), .Q(
        \RegFilePlugin_regFile[4][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][11]  ( .D(n4311), .CP(n7247), .Q(
        \RegFilePlugin_regFile[3][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][11]  ( .D(n4279), .CP(n7151), .Q(
        \RegFilePlugin_regFile[2][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][11]  ( .D(n4247), .CP(n7247), .Q(
        \RegFilePlugin_regFile[1][11] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][11]  ( .D(n4174), .CP(n7247), .Q(
        \RegFilePlugin_regFile[0][11] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[11]  ( .D(N843), .CP(n7153), .Q(
        _zz_RegFilePlugin_regFile_port0[11]) );
  dfnrq1 \decode_to_execute_RS1_reg[11]  ( .D(n4173), .CP(n7155), .Q(
        execute_RS1[11]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[11]  ( .D(n6144), .CP(
        n7158), .Q(_zz_CsrPlugin_csrMapping_readDataInit[11]) );
  dfnrq1 CsrPlugin_mie_MEIE_reg ( .D(n6130), .CP(n7159), .Q(CsrPlugin_mie_MEIE) );
  dfnrq1 \CsrPlugin_mstatus_MPP_reg[0]  ( .D(n6127), .CP(n7153), .Q(
        CsrPlugin_mstatus_MPP[0]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[9]  ( .D(n4132), .CP(n7155), .Q(
        CsrPlugin_mtvec_base[9]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[11]  ( .D(n6108), .CP(n7157), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[11]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[11]  ( .D(n5895), .CP(
        n7157), .Q(iBusWishbone_ADR[9]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[11]  ( 
        .D(n5258), .CP(n7157), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[11]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[11]  ( .D(
        n6186), .CP(n7157), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[11]) );
  dfnrq1 \CsrPlugin_mtval_reg[11]  ( .D(n6018), .CP(n7157), .Q(
        CsrPlugin_mtval[11]) );
  dfnrq1 \decode_to_execute_PC_reg[11]  ( .D(n5257), .CP(n7157), .Q(
        execute_PC[11]) );
  dfnrq1 \memory_to_writeBack_PC_reg[11]  ( .D(n5256), .CP(n7157), .Q(
        writeBack_PC[11]) );
  dfnrq1 \CsrPlugin_mepc_reg[11]  ( .D(n4100), .CP(n7157), .Q(
        CsrPlugin_mepc[11]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[11]  ( .D(n6061), .CP(n7156), .Q(
        debug_bus_rsp_data[11]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[11]  ( .D(N876), .CP(n7156), .Q(
        _zz_RegFilePlugin_regFile_port1[11]) );
  dfnrq1 \decode_to_execute_RS2_reg[11]  ( .D(n4172), .CP(n7156), .Q(
        execute_RS2[11]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][10]  ( .D(n5206), .CP(n7156), .Q(
        \RegFilePlugin_regFile[31][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][10]  ( .D(n5174), .CP(n7156), .Q(
        \RegFilePlugin_regFile[30][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][10]  ( .D(n5142), .CP(n7156), .Q(
        \RegFilePlugin_regFile[29][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][10]  ( .D(n5110), .CP(n7156), .Q(
        \RegFilePlugin_regFile[28][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][10]  ( .D(n5078), .CP(n7156), .Q(
        \RegFilePlugin_regFile[27][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][10]  ( .D(n5046), .CP(n7155), .Q(
        \RegFilePlugin_regFile[26][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][10]  ( .D(n5014), .CP(n7155), .Q(
        \RegFilePlugin_regFile[25][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][10]  ( .D(n4982), .CP(n7155), .Q(
        \RegFilePlugin_regFile[24][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][10]  ( .D(n4950), .CP(n7155), .Q(
        \RegFilePlugin_regFile[23][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][10]  ( .D(n4918), .CP(n7155), .Q(
        \RegFilePlugin_regFile[22][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][10]  ( .D(n4886), .CP(n7155), .Q(
        \RegFilePlugin_regFile[21][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][10]  ( .D(n4854), .CP(n7155), .Q(
        \RegFilePlugin_regFile[20][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][10]  ( .D(n4822), .CP(n7155), .Q(
        \RegFilePlugin_regFile[19][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][10]  ( .D(n4790), .CP(n7159), .Q(
        \RegFilePlugin_regFile[18][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][10]  ( .D(n4758), .CP(n7152), .Q(
        \RegFilePlugin_regFile[17][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][10]  ( .D(n4726), .CP(n7156), .Q(
        \RegFilePlugin_regFile[16][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][10]  ( .D(n4694), .CP(n7260), .Q(
        \RegFilePlugin_regFile[15][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][10]  ( .D(n4662), .CP(n7246), .Q(
        \RegFilePlugin_regFile[14][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][10]  ( .D(n4630), .CP(n7158), .Q(
        \RegFilePlugin_regFile[13][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][10]  ( .D(n4598), .CP(n7157), .Q(
        \RegFilePlugin_regFile[12][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][10]  ( .D(n4566), .CP(n7151), .Q(
        \RegFilePlugin_regFile[11][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][10]  ( .D(n4534), .CP(n7154), .Q(
        \RegFilePlugin_regFile[10][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][10]  ( .D(n4502), .CP(n7154), .Q(
        \RegFilePlugin_regFile[9][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][10]  ( .D(n4470), .CP(n7154), .Q(
        \RegFilePlugin_regFile[8][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][10]  ( .D(n4438), .CP(n7154), .Q(
        \RegFilePlugin_regFile[7][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][10]  ( .D(n4406), .CP(n7154), .Q(
        \RegFilePlugin_regFile[6][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][10]  ( .D(n4374), .CP(n7154), .Q(
        \RegFilePlugin_regFile[5][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][10]  ( .D(n4342), .CP(n7154), .Q(
        \RegFilePlugin_regFile[4][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][10]  ( .D(n4310), .CP(n7154), .Q(
        \RegFilePlugin_regFile[3][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][10]  ( .D(n4278), .CP(n7246), .Q(
        \RegFilePlugin_regFile[2][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][10]  ( .D(n4246), .CP(n7156), .Q(
        \RegFilePlugin_regFile[1][10] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][10]  ( .D(n4171), .CP(n7152), .Q(
        \RegFilePlugin_regFile[0][10] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[10]  ( .D(N844), .CP(n7152), .Q(
        _zz_RegFilePlugin_regFile_port0[10]) );
  dfnrq1 \decode_to_execute_RS1_reg[10]  ( .D(n4170), .CP(n7151), .Q(
        execute_RS1[10]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[10]  ( .D(n6143), .CP(
        n7158), .Q(_zz_CsrPlugin_csrMapping_readDataInit[10]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[8]  ( .D(n4133), .CP(n7157), .Q(
        CsrPlugin_mtvec_base[8]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[10]  ( .D(n6109), .CP(n7153), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[10]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[10]  ( .D(n5894), .CP(
        n7159), .Q(iBusWishbone_ADR[8]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[10]  ( 
        .D(n5255), .CP(n7156), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[10]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[10]  ( .D(
        n6185), .CP(n7260), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[10]) );
  dfnrq1 \CsrPlugin_mtval_reg[10]  ( .D(n6017), .CP(n7152), .Q(
        CsrPlugin_mtval[10]) );
  dfnrq1 \decode_to_execute_PC_reg[10]  ( .D(n5254), .CP(n7151), .Q(
        execute_PC[10]) );
  dfnrq1 \memory_to_writeBack_PC_reg[10]  ( .D(n5253), .CP(n7158), .Q(
        writeBack_PC[10]) );
  dfnrq1 \CsrPlugin_mepc_reg[10]  ( .D(n4101), .CP(n7157), .Q(
        CsrPlugin_mepc[10]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[10]  ( .D(n6062), .CP(n7153), .Q(
        debug_bus_rsp_data[10]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[10]  ( .D(N877), .CP(n7154), .Q(
        _zz_RegFilePlugin_regFile_port1[10]) );
  dfnrq1 \decode_to_execute_RS2_reg[10]  ( .D(n4169), .CP(n7157), .Q(
        execute_RS2[10]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][9]  ( .D(n5205), .CP(n7158), .Q(
        \RegFilePlugin_regFile[31][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][9]  ( .D(n5173), .CP(n7151), .Q(
        \RegFilePlugin_regFile[30][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][9]  ( .D(n5141), .CP(n7152), .Q(
        \RegFilePlugin_regFile[29][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][9]  ( .D(n5109), .CP(n7156), .Q(
        \RegFilePlugin_regFile[28][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][9]  ( .D(n5077), .CP(n7247), .Q(
        \RegFilePlugin_regFile[27][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][9]  ( .D(n5045), .CP(n7157), .Q(
        \RegFilePlugin_regFile[26][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][9]  ( .D(n5013), .CP(n7153), .Q(
        \RegFilePlugin_regFile[25][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][9]  ( .D(n4981), .CP(n7153), .Q(
        \RegFilePlugin_regFile[24][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][9]  ( .D(n4949), .CP(n7153), .Q(
        \RegFilePlugin_regFile[23][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][9]  ( .D(n4917), .CP(n7153), .Q(
        \RegFilePlugin_regFile[22][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][9]  ( .D(n4885), .CP(n7153), .Q(
        \RegFilePlugin_regFile[21][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][9]  ( .D(n4853), .CP(n7153), .Q(
        \RegFilePlugin_regFile[20][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][9]  ( .D(n4821), .CP(n7153), .Q(
        \RegFilePlugin_regFile[19][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][9]  ( .D(n4789), .CP(n7153), .Q(
        \RegFilePlugin_regFile[18][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][9]  ( .D(n4757), .CP(n7152), .Q(
        \RegFilePlugin_regFile[17][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][9]  ( .D(n4725), .CP(n7152), .Q(
        \RegFilePlugin_regFile[16][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][9]  ( .D(n4693), .CP(n7152), .Q(
        \RegFilePlugin_regFile[15][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][9]  ( .D(n4661), .CP(n7152), .Q(
        \RegFilePlugin_regFile[14][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][9]  ( .D(n4629), .CP(n7152), .Q(
        \RegFilePlugin_regFile[13][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][9]  ( .D(n4597), .CP(n7152), .Q(
        \RegFilePlugin_regFile[12][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][9]  ( .D(n4565), .CP(n7152), .Q(
        \RegFilePlugin_regFile[11][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][9]  ( .D(n4533), .CP(n7152), .Q(
        \RegFilePlugin_regFile[10][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][9]  ( .D(n4501), .CP(n7151), .Q(
        \RegFilePlugin_regFile[9][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][9]  ( .D(n4469), .CP(n7154), .Q(
        \RegFilePlugin_regFile[8][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][9]  ( .D(n4437), .CP(n7158), .Q(
        \RegFilePlugin_regFile[7][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][9]  ( .D(n4405), .CP(n7154), .Q(
        \RegFilePlugin_regFile[6][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][9]  ( .D(n4373), .CP(n7157), .Q(
        \RegFilePlugin_regFile[5][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][9]  ( .D(n4341), .CP(n7154), .Q(
        \RegFilePlugin_regFile[4][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][9]  ( .D(n4309), .CP(n7153), .Q(
        \RegFilePlugin_regFile[3][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][9]  ( .D(n4277), .CP(n7154), .Q(
        \RegFilePlugin_regFile[2][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][9]  ( .D(n4245), .CP(n7151), .Q(
        \RegFilePlugin_regFile[1][9] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][9]  ( .D(n4168), .CP(n7151), .Q(
        \RegFilePlugin_regFile[0][9] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[9]  ( .D(N845), .CP(n7151), .Q(
        _zz_RegFilePlugin_regFile_port0[9]) );
  dfnrq1 \decode_to_execute_RS1_reg[9]  ( .D(n4167), .CP(n7151), .Q(
        execute_RS1[9]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[9]  ( .D(n6142), .CP(n7151), .Q(_zz_CsrPlugin_csrMapping_readDataInit[9]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[7]  ( .D(n4134), .CP(n7151), .Q(
        CsrPlugin_mtvec_base[7]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[9]  ( .D(n6110), .CP(n7151), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[9]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[9]  ( .D(n5893), .CP(
        n7151), .Q(iBusWishbone_ADR[7]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[9]  ( 
        .D(n5252), .CP(n7142), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[9]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[9]  ( .D(
        n6184), .CP(n7149), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[9]) );
  dfnrq1 \CsrPlugin_mtval_reg[9]  ( .D(n6016), .CP(n7148), .Q(
        CsrPlugin_mtval[9]) );
  dfnrq1 \decode_to_execute_PC_reg[9]  ( .D(n5251), .CP(n7144), .Q(
        execute_PC[9]) );
  dfnrq1 \memory_to_writeBack_PC_reg[9]  ( .D(n5250), .CP(n7146), .Q(
        writeBack_PC[9]) );
  dfnrq1 \CsrPlugin_mepc_reg[9]  ( .D(n4102), .CP(n7249), .Q(CsrPlugin_mepc[9]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[9]  ( .D(n6063), .CP(n7150), .Q(
        debug_bus_rsp_data[9]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[9]  ( .D(N878), .CP(n7248), .Q(
        _zz_RegFilePlugin_regFile_port1[9]) );
  dfnrq1 \decode_to_execute_RS2_reg[9]  ( .D(n4166), .CP(n7148), .Q(
        execute_RS2[9]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][8]  ( .D(n5204), .CP(n7149), .Q(
        \RegFilePlugin_regFile[31][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][8]  ( .D(n5172), .CP(n7261), .Q(
        \RegFilePlugin_regFile[30][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][8]  ( .D(n5140), .CP(n7248), .Q(
        \RegFilePlugin_regFile[29][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][8]  ( .D(n5108), .CP(n7147), .Q(
        \RegFilePlugin_regFile[28][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][8]  ( .D(n5076), .CP(n7147), .Q(
        \RegFilePlugin_regFile[27][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][8]  ( .D(n5044), .CP(n7143), .Q(
        \RegFilePlugin_regFile[26][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][8]  ( .D(n5012), .CP(n7142), .Q(
        \RegFilePlugin_regFile[25][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][8]  ( .D(n4980), .CP(n7261), .Q(
        \RegFilePlugin_regFile[24][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][8]  ( .D(n4948), .CP(n7149), .Q(
        \RegFilePlugin_regFile[23][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][8]  ( .D(n4916), .CP(n7148), .Q(
        \RegFilePlugin_regFile[22][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][8]  ( .D(n4884), .CP(n7261), .Q(
        \RegFilePlugin_regFile[21][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][8]  ( .D(n4852), .CP(n7149), .Q(
        \RegFilePlugin_regFile[20][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][8]  ( .D(n4820), .CP(n7261), .Q(
        \RegFilePlugin_regFile[19][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][8]  ( .D(n4788), .CP(n7248), .Q(
        \RegFilePlugin_regFile[18][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][8]  ( .D(n4756), .CP(n7147), .Q(
        \RegFilePlugin_regFile[17][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][8]  ( .D(n4724), .CP(n7147), .Q(
        \RegFilePlugin_regFile[16][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][8]  ( .D(n4692), .CP(n7143), .Q(
        \RegFilePlugin_regFile[15][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][8]  ( .D(n4660), .CP(n7248), .Q(
        \RegFilePlugin_regFile[14][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][8]  ( .D(n4628), .CP(n7146), .Q(
        \RegFilePlugin_regFile[13][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][8]  ( .D(n4596), .CP(n7142), .Q(
        \RegFilePlugin_regFile[12][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][8]  ( .D(n4564), .CP(n7261), .Q(
        \RegFilePlugin_regFile[11][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][8]  ( .D(n4532), .CP(n7143), .Q(
        \RegFilePlugin_regFile[10][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][8]  ( .D(n4500), .CP(n7145), .Q(
        \RegFilePlugin_regFile[9][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][8]  ( .D(n4468), .CP(n7248), .Q(
        \RegFilePlugin_regFile[8][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][8]  ( .D(n4436), .CP(n7248), .Q(
        \RegFilePlugin_regFile[7][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][8]  ( .D(n4404), .CP(n7248), .Q(
        \RegFilePlugin_regFile[6][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][8]  ( .D(n4372), .CP(n7248), .Q(
        \RegFilePlugin_regFile[5][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][8]  ( .D(n4340), .CP(n7145), .Q(
        \RegFilePlugin_regFile[4][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][8]  ( .D(n4308), .CP(n7149), .Q(
        \RegFilePlugin_regFile[3][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][8]  ( .D(n4276), .CP(n7248), .Q(
        \RegFilePlugin_regFile[2][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][8]  ( .D(n4244), .CP(n7142), .Q(
        \RegFilePlugin_regFile[1][8] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][8]  ( .D(n4165), .CP(n7248), .Q(
        \RegFilePlugin_regFile[0][8] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[8]  ( .D(N846), .CP(n7248), .Q(
        _zz_RegFilePlugin_regFile_port0[8]) );
  dfnrq1 \decode_to_execute_RS1_reg[8]  ( .D(n4164), .CP(n7145), .Q(
        execute_RS1[8]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[8]  ( .D(n6141), .CP(n7143), .Q(_zz_CsrPlugin_csrMapping_readDataInit[8]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[6]  ( .D(n4135), .CP(n7248), .Q(
        CsrPlugin_mtvec_base[6]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[8]  ( .D(n6111), .CP(n7145), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[8]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[8]  ( .D(n5892), .CP(
        n7143), .Q(iBusWishbone_ADR[6]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[8]  ( 
        .D(n5249), .CP(n7142), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[8]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[8]  ( .D(
        n6183), .CP(n7150), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[8]) );
  dfnrq1 \CsrPlugin_mtval_reg[8]  ( .D(n6015), .CP(n7150), .Q(
        CsrPlugin_mtval[8]) );
  dfnrq1 \decode_to_execute_PC_reg[8]  ( .D(n5248), .CP(n7150), .Q(
        execute_PC[8]) );
  dfnrq1 \memory_to_writeBack_PC_reg[8]  ( .D(n5247), .CP(n7150), .Q(
        writeBack_PC[8]) );
  dfnrq1 \CsrPlugin_mepc_reg[8]  ( .D(n4103), .CP(n7150), .Q(CsrPlugin_mepc[8]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[8]  ( .D(n6064), .CP(n7150), .Q(
        debug_bus_rsp_data[8]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[8]  ( .D(N879), .CP(n7150), .Q(
        _zz_RegFilePlugin_regFile_port1[8]) );
  dfnrq1 \decode_to_execute_RS2_reg[8]  ( .D(n4163), .CP(n7150), .Q(
        execute_RS2[8]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][7]  ( .D(n5203), .CP(n7149), .Q(
        \RegFilePlugin_regFile[31][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][7]  ( .D(n5171), .CP(n7149), .Q(
        \RegFilePlugin_regFile[30][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][7]  ( .D(n5139), .CP(n7149), .Q(
        \RegFilePlugin_regFile[29][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][7]  ( .D(n5107), .CP(n7149), .Q(
        \RegFilePlugin_regFile[28][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][7]  ( .D(n5075), .CP(n7149), .Q(
        \RegFilePlugin_regFile[27][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][7]  ( .D(n5043), .CP(n7149), .Q(
        \RegFilePlugin_regFile[26][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][7]  ( .D(n5011), .CP(n7149), .Q(
        \RegFilePlugin_regFile[25][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][7]  ( .D(n4979), .CP(n7149), .Q(
        \RegFilePlugin_regFile[24][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][7]  ( .D(n4947), .CP(n7146), .Q(
        \RegFilePlugin_regFile[23][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][7]  ( .D(n4915), .CP(n7146), .Q(
        \RegFilePlugin_regFile[22][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][7]  ( .D(n4883), .CP(n7146), .Q(
        \RegFilePlugin_regFile[21][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][7]  ( .D(n4851), .CP(n7249), .Q(
        \RegFilePlugin_regFile[20][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][7]  ( .D(n4819), .CP(n7146), .Q(
        \RegFilePlugin_regFile[19][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][7]  ( .D(n4787), .CP(n7249), .Q(
        \RegFilePlugin_regFile[18][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][7]  ( .D(n4755), .CP(n7146), .Q(
        \RegFilePlugin_regFile[17][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][7]  ( .D(n4723), .CP(n7249), .Q(
        \RegFilePlugin_regFile[16][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][7]  ( .D(n4691), .CP(n7144), .Q(
        \RegFilePlugin_regFile[15][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][7]  ( .D(n4659), .CP(n7144), .Q(
        \RegFilePlugin_regFile[14][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][7]  ( .D(n4627), .CP(n7144), .Q(
        \RegFilePlugin_regFile[13][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][7]  ( .D(n4595), .CP(n7150), .Q(
        \RegFilePlugin_regFile[12][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][7]  ( .D(n4563), .CP(n7144), .Q(
        \RegFilePlugin_regFile[11][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][7]  ( .D(n4531), .CP(n7150), .Q(
        \RegFilePlugin_regFile[10][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][7]  ( .D(n4499), .CP(n7144), .Q(
        \RegFilePlugin_regFile[9][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][7]  ( .D(n4467), .CP(n7150), .Q(
        \RegFilePlugin_regFile[8][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][7]  ( .D(n4435), .CP(n7261), .Q(
        \RegFilePlugin_regFile[7][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][7]  ( .D(n4403), .CP(n7148), .Q(
        \RegFilePlugin_regFile[6][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][7]  ( .D(n4371), .CP(n7261), .Q(
        \RegFilePlugin_regFile[5][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][7]  ( .D(n4339), .CP(n7249), .Q(
        \RegFilePlugin_regFile[4][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][7]  ( .D(n4307), .CP(n7261), .Q(
        \RegFilePlugin_regFile[3][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][7]  ( .D(n4275), .CP(n7261), .Q(
        \RegFilePlugin_regFile[2][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][7]  ( .D(n4243), .CP(n7261), .Q(
        \RegFilePlugin_regFile[1][7] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][7]  ( .D(n4162), .CP(n7150), .Q(
        \RegFilePlugin_regFile[0][7] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[7]  ( .D(N847), .CP(n7261), .Q(
        _zz_RegFilePlugin_regFile_port0[7]) );
  dfnrq1 \decode_to_execute_RS1_reg[7]  ( .D(n4161), .CP(n7261), .Q(
        execute_RS1[7]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[7]  ( .D(n6140), .CP(n7261), .Q(_zz_CsrPlugin_csrMapping_readDataInit[7]) );
  dfnrq1 CsrPlugin_mie_MTIE_reg ( .D(n6128), .CP(n7261), .Q(CsrPlugin_mie_MTIE) );
  dfnrq1 CsrPlugin_mstatus_MPIE_reg ( .D(n6125), .CP(n7146), .Q(
        CsrPlugin_mstatus_MPIE) );
  dfnrq1 CsrPlugin_mstatus_MIE_reg ( .D(n6124), .CP(n7249), .Q(
        CsrPlugin_mstatus_MIE) );
  dfnrq1 CsrPlugin_interrupt_valid_reg ( .D(N1785), .CP(n7261), .Q(
        CsrPlugin_interrupt_valid) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[5]  ( .D(n4136), .CP(n7261), .Q(
        CsrPlugin_mtvec_base[5]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[7]  ( .D(n6112), .CP(n7249), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[7]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[7]  ( .D(n5891), .CP(
        n7249), .Q(iBusWishbone_ADR[5]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[7]  ( 
        .D(n5246), .CP(n7147), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[7]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[7]  ( .D(
        n6182), .CP(n7249), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[7]) );
  dfnrq1 \CsrPlugin_mtval_reg[7]  ( .D(n6014), .CP(n7147), .Q(
        CsrPlugin_mtval[7]) );
  dfnrq1 \decode_to_execute_PC_reg[7]  ( .D(n5245), .CP(n7248), .Q(
        execute_PC[7]) );
  dfnrq1 \memory_to_writeBack_PC_reg[7]  ( .D(n5244), .CP(n7148), .Q(
        writeBack_PC[7]) );
  dfnrq1 \CsrPlugin_mepc_reg[7]  ( .D(n4104), .CP(n7249), .Q(CsrPlugin_mepc[7]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[7]  ( .D(n6065), .CP(n7249), .Q(
        debug_bus_rsp_data[7]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[7]  ( .D(N880), .CP(n7248), .Q(
        _zz_RegFilePlugin_regFile_port1[7]) );
  dfnrq1 \decode_to_execute_RS2_reg[7]  ( .D(n4160), .CP(n7150), .Q(
        execute_RS2[7]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][6]  ( .D(n5202), .CP(n7143), .Q(
        \RegFilePlugin_regFile[31][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][6]  ( .D(n5170), .CP(n7249), .Q(
        \RegFilePlugin_regFile[30][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][6]  ( .D(n5138), .CP(n7248), .Q(
        \RegFilePlugin_regFile[29][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][6]  ( .D(n5106), .CP(n7249), .Q(
        \RegFilePlugin_regFile[28][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][6]  ( .D(n5074), .CP(n7142), .Q(
        \RegFilePlugin_regFile[27][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][6]  ( .D(n5042), .CP(n7249), .Q(
        \RegFilePlugin_regFile[26][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][6]  ( .D(n5010), .CP(n7249), .Q(
        \RegFilePlugin_regFile[25][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][6]  ( .D(n4978), .CP(n7144), .Q(
        \RegFilePlugin_regFile[24][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][6]  ( .D(n4946), .CP(n7146), .Q(
        \RegFilePlugin_regFile[23][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][6]  ( .D(n4914), .CP(n7149), .Q(
        \RegFilePlugin_regFile[22][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][6]  ( .D(n4882), .CP(n7150), .Q(
        \RegFilePlugin_regFile[21][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][6]  ( .D(n4850), .CP(n7144), .Q(
        \RegFilePlugin_regFile[20][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][6]  ( .D(n4818), .CP(n7146), .Q(
        \RegFilePlugin_regFile[19][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][6]  ( .D(n4786), .CP(n7148), .Q(
        \RegFilePlugin_regFile[18][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][6]  ( .D(n4754), .CP(n7148), .Q(
        \RegFilePlugin_regFile[17][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][6]  ( .D(n4722), .CP(n7148), .Q(
        \RegFilePlugin_regFile[16][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][6]  ( .D(n4690), .CP(n7148), .Q(
        \RegFilePlugin_regFile[15][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][6]  ( .D(n4658), .CP(n7148), .Q(
        \RegFilePlugin_regFile[14][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][6]  ( .D(n4626), .CP(n7148), .Q(
        \RegFilePlugin_regFile[13][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][6]  ( .D(n4594), .CP(n7148), .Q(
        \RegFilePlugin_regFile[12][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][6]  ( .D(n4562), .CP(n7148), .Q(
        \RegFilePlugin_regFile[11][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][6]  ( .D(n4530), .CP(n7147), .Q(
        \RegFilePlugin_regFile[10][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][6]  ( .D(n4498), .CP(n7147), .Q(
        \RegFilePlugin_regFile[9][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][6]  ( .D(n4466), .CP(n7147), .Q(
        \RegFilePlugin_regFile[8][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][6]  ( .D(n4434), .CP(n7147), .Q(
        \RegFilePlugin_regFile[7][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][6]  ( .D(n4402), .CP(n7147), .Q(
        \RegFilePlugin_regFile[6][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][6]  ( .D(n4370), .CP(n7147), .Q(
        \RegFilePlugin_regFile[5][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][6]  ( .D(n4338), .CP(n7147), .Q(
        \RegFilePlugin_regFile[4][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][6]  ( .D(n4306), .CP(n7147), .Q(
        \RegFilePlugin_regFile[3][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][6]  ( .D(n4274), .CP(n7146), .Q(
        \RegFilePlugin_regFile[2][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][6]  ( .D(n4242), .CP(n7146), .Q(
        \RegFilePlugin_regFile[1][6] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][6]  ( .D(n4159), .CP(n7146), .Q(
        \RegFilePlugin_regFile[0][6] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[6]  ( .D(N848), .CP(n7146), .Q(
        _zz_RegFilePlugin_regFile_port0[6]) );
  dfnrq1 \decode_to_execute_RS1_reg[6]  ( .D(n4158), .CP(n7146), .Q(
        execute_RS1[6]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[6]  ( .D(n6139), .CP(n7146), .Q(_zz_CsrPlugin_csrMapping_readDataInit[6]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[4]  ( .D(n4137), .CP(n7146), .Q(
        CsrPlugin_mtvec_base[4]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[6]  ( .D(n6113), .CP(n7146), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[6]) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_address_reg[6]  ( .D(n5890), .CP(
        n7150), .Q(iBusWishbone_ADR[4]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[6]  ( 
        .D(n5243), .CP(n7143), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[6]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[6]  ( .D(
        n6181), .CP(n7147), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[6]) );
  dfnrq1 \CsrPlugin_mtval_reg[6]  ( .D(n6013), .CP(n7261), .Q(
        CsrPlugin_mtval[6]) );
  dfnrq1 \decode_to_execute_PC_reg[6]  ( .D(n5242), .CP(n7248), .Q(
        execute_PC[6]) );
  dfnrq1 \memory_to_writeBack_PC_reg[6]  ( .D(n5241), .CP(n7149), .Q(
        writeBack_PC[6]) );
  dfnrq1 \CsrPlugin_mepc_reg[6]  ( .D(n4105), .CP(n7148), .Q(CsrPlugin_mepc[6]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[6]  ( .D(n6066), .CP(n7142), .Q(
        debug_bus_rsp_data[6]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[6]  ( .D(N881), .CP(n7145), .Q(
        _zz_RegFilePlugin_regFile_port1[6]) );
  dfnrq1 \decode_to_execute_RS2_reg[6]  ( .D(n4157), .CP(n7145), .Q(
        execute_RS2[6]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][5]  ( .D(n5201), .CP(n7145), .Q(
        \RegFilePlugin_regFile[31][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][5]  ( .D(n5169), .CP(n7145), .Q(
        \RegFilePlugin_regFile[30][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][5]  ( .D(n5137), .CP(n7145), .Q(
        \RegFilePlugin_regFile[29][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][5]  ( .D(n5105), .CP(n7145), .Q(
        \RegFilePlugin_regFile[28][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][5]  ( .D(n5073), .CP(n7145), .Q(
        \RegFilePlugin_regFile[27][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][5]  ( .D(n5041), .CP(n7145), .Q(
        \RegFilePlugin_regFile[26][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][5]  ( .D(n5009), .CP(n7248), .Q(
        \RegFilePlugin_regFile[25][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][5]  ( .D(n4977), .CP(n7147), .Q(
        \RegFilePlugin_regFile[24][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][5]  ( .D(n4945), .CP(n7143), .Q(
        \RegFilePlugin_regFile[23][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][5]  ( .D(n4913), .CP(n7143), .Q(
        \RegFilePlugin_regFile[22][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][5]  ( .D(n4881), .CP(n7142), .Q(
        \RegFilePlugin_regFile[21][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][5]  ( .D(n4849), .CP(n7149), .Q(
        \RegFilePlugin_regFile[20][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][5]  ( .D(n4817), .CP(n7148), .Q(
        \RegFilePlugin_regFile[19][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][5]  ( .D(n4785), .CP(n7144), .Q(
        \RegFilePlugin_regFile[18][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][5]  ( .D(n4753), .CP(n7150), .Q(
        \RegFilePlugin_regFile[17][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][5]  ( .D(n4721), .CP(n7147), .Q(
        \RegFilePlugin_regFile[16][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][5]  ( .D(n4689), .CP(n7261), .Q(
        \RegFilePlugin_regFile[15][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][5]  ( .D(n4657), .CP(n7143), .Q(
        \RegFilePlugin_regFile[14][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][5]  ( .D(n4625), .CP(n7142), .Q(
        \RegFilePlugin_regFile[13][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][5]  ( .D(n4593), .CP(n7149), .Q(
        \RegFilePlugin_regFile[12][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][5]  ( .D(n4561), .CP(n7148), .Q(
        \RegFilePlugin_regFile[11][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][5]  ( .D(n4529), .CP(n7144), .Q(
        \RegFilePlugin_regFile[10][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][5]  ( .D(n4497), .CP(n7145), .Q(
        \RegFilePlugin_regFile[9][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][5]  ( .D(n4465), .CP(n7148), .Q(
        \RegFilePlugin_regFile[8][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][5]  ( .D(n4433), .CP(n7149), .Q(
        \RegFilePlugin_regFile[7][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][5]  ( .D(n4401), .CP(n7142), .Q(
        \RegFilePlugin_regFile[6][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][5]  ( .D(n4369), .CP(n7143), .Q(
        \RegFilePlugin_regFile[5][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][5]  ( .D(n4337), .CP(n7147), .Q(
        \RegFilePlugin_regFile[4][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][5]  ( .D(n4305), .CP(n7249), .Q(
        \RegFilePlugin_regFile[3][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][5]  ( .D(n4273), .CP(n7148), .Q(
        \RegFilePlugin_regFile[2][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][5]  ( .D(n4241), .CP(n7144), .Q(
        \RegFilePlugin_regFile[1][5] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][5]  ( .D(n4156), .CP(n7144), .Q(
        \RegFilePlugin_regFile[0][5] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[5]  ( .D(N849), .CP(n7144), .Q(
        _zz_RegFilePlugin_regFile_port0[5]) );
  dfnrq1 \decode_to_execute_RS1_reg[5]  ( .D(n4155), .CP(n7144), .Q(
        execute_RS1[5]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[5]  ( .D(N882), .CP(n7144), .Q(
        _zz_RegFilePlugin_regFile_port1[5]) );
  dfnrq1 \decode_to_execute_RS2_reg[5]  ( .D(n4154), .CP(n7144), .Q(
        execute_RS2[5]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][4]  ( .D(n5200), .CP(n7144), .Q(
        \RegFilePlugin_regFile[31][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][4]  ( .D(n5168), .CP(n7144), .Q(
        \RegFilePlugin_regFile[30][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][4]  ( .D(n5136), .CP(n7143), .Q(
        \RegFilePlugin_regFile[29][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][4]  ( .D(n5104), .CP(n7143), .Q(
        \RegFilePlugin_regFile[28][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][4]  ( .D(n5072), .CP(n7143), .Q(
        \RegFilePlugin_regFile[27][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][4]  ( .D(n5040), .CP(n7143), .Q(
        \RegFilePlugin_regFile[26][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][4]  ( .D(n5008), .CP(n7143), .Q(
        \RegFilePlugin_regFile[25][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][4]  ( .D(n4976), .CP(n7143), .Q(
        \RegFilePlugin_regFile[24][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][4]  ( .D(n4944), .CP(n7143), .Q(
        \RegFilePlugin_regFile[23][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][4]  ( .D(n4912), .CP(n7143), .Q(
        \RegFilePlugin_regFile[22][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][4]  ( .D(n4880), .CP(n7142), .Q(
        \RegFilePlugin_regFile[21][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][4]  ( .D(n4848), .CP(n7145), .Q(
        \RegFilePlugin_regFile[20][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][4]  ( .D(n4816), .CP(n7149), .Q(
        \RegFilePlugin_regFile[19][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][4]  ( .D(n4784), .CP(n7145), .Q(
        \RegFilePlugin_regFile[18][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][4]  ( .D(n4752), .CP(n7148), .Q(
        \RegFilePlugin_regFile[17][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][4]  ( .D(n4720), .CP(n7145), .Q(
        \RegFilePlugin_regFile[16][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][4]  ( .D(n4688), .CP(n7144), .Q(
        \RegFilePlugin_regFile[15][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][4]  ( .D(n4656), .CP(n7145), .Q(
        \RegFilePlugin_regFile[14][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][4]  ( .D(n4624), .CP(n7142), .Q(
        \RegFilePlugin_regFile[13][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][4]  ( .D(n4592), .CP(n7142), .Q(
        \RegFilePlugin_regFile[12][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][4]  ( .D(n4560), .CP(n7142), .Q(
        \RegFilePlugin_regFile[11][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][4]  ( .D(n4528), .CP(n7142), .Q(
        \RegFilePlugin_regFile[10][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][4]  ( .D(n4496), .CP(n7142), .Q(
        \RegFilePlugin_regFile[9][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][4]  ( .D(n4464), .CP(n7142), .Q(
        \RegFilePlugin_regFile[8][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][4]  ( .D(n4432), .CP(n7142), .Q(
        \RegFilePlugin_regFile[7][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][4]  ( .D(n4400), .CP(n7142), .Q(
        \RegFilePlugin_regFile[6][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][4]  ( .D(n4368), .CP(n7133), .Q(
        \RegFilePlugin_regFile[5][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][4]  ( .D(n4336), .CP(n7140), .Q(
        \RegFilePlugin_regFile[4][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][4]  ( .D(n4304), .CP(n7139), .Q(
        \RegFilePlugin_regFile[3][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][4]  ( .D(n4272), .CP(n7135), .Q(
        \RegFilePlugin_regFile[2][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][4]  ( .D(n4240), .CP(n7137), .Q(
        \RegFilePlugin_regFile[1][4] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][4]  ( .D(n4153), .CP(n7251), .Q(
        \RegFilePlugin_regFile[0][4] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[4]  ( .D(N850), .CP(n7141), .Q(
        _zz_RegFilePlugin_regFile_port0[4]) );
  dfnrq1 \decode_to_execute_RS1_reg[4]  ( .D(n4152), .CP(n7250), .Q(
        execute_RS1[4]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[4]  ( .D(N883), .CP(n7139), .Q(
        _zz_RegFilePlugin_regFile_port1[4]) );
  dfnrq1 \decode_to_execute_RS2_reg[4]  ( .D(n4151), .CP(n7140), .Q(
        execute_RS2[4]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[3]  ( .D(n6069), .CP(n7262), .Q(
        DebugPlugin_busReadDataReg[3]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][3]  ( .D(n5199), .CP(n7250), .Q(
        \RegFilePlugin_regFile[31][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][3]  ( .D(n5167), .CP(n7138), .Q(
        \RegFilePlugin_regFile[30][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][3]  ( .D(n5135), .CP(n7138), .Q(
        \RegFilePlugin_regFile[29][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][3]  ( .D(n5103), .CP(n7134), .Q(
        \RegFilePlugin_regFile[28][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][3]  ( .D(n5071), .CP(n7133), .Q(
        \RegFilePlugin_regFile[27][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][3]  ( .D(n5039), .CP(n7262), .Q(
        \RegFilePlugin_regFile[26][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][3]  ( .D(n5007), .CP(n7140), .Q(
        \RegFilePlugin_regFile[25][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][3]  ( .D(n4975), .CP(n7139), .Q(
        \RegFilePlugin_regFile[24][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][3]  ( .D(n4943), .CP(n7262), .Q(
        \RegFilePlugin_regFile[23][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][3]  ( .D(n4911), .CP(n7140), .Q(
        \RegFilePlugin_regFile[22][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][3]  ( .D(n4879), .CP(n7262), .Q(
        \RegFilePlugin_regFile[21][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][3]  ( .D(n4847), .CP(n7250), .Q(
        \RegFilePlugin_regFile[20][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][3]  ( .D(n4815), .CP(n7138), .Q(
        \RegFilePlugin_regFile[19][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][3]  ( .D(n4783), .CP(n7138), .Q(
        \RegFilePlugin_regFile[18][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][3]  ( .D(n4751), .CP(n7134), .Q(
        \RegFilePlugin_regFile[17][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][3]  ( .D(n4719), .CP(n7250), .Q(
        \RegFilePlugin_regFile[16][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][3]  ( .D(n4687), .CP(n7137), .Q(
        \RegFilePlugin_regFile[15][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][3]  ( .D(n4655), .CP(n7133), .Q(
        \RegFilePlugin_regFile[14][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][3]  ( .D(n4623), .CP(n7262), .Q(
        \RegFilePlugin_regFile[13][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][3]  ( .D(n4591), .CP(n7134), .Q(
        \RegFilePlugin_regFile[12][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][3]  ( .D(n4559), .CP(n7136), .Q(
        \RegFilePlugin_regFile[11][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][3]  ( .D(n4527), .CP(n7250), .Q(
        \RegFilePlugin_regFile[10][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][3]  ( .D(n4495), .CP(n7250), .Q(
        \RegFilePlugin_regFile[9][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][3]  ( .D(n4463), .CP(n7250), .Q(
        \RegFilePlugin_regFile[8][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][3]  ( .D(n4431), .CP(n7250), .Q(
        \RegFilePlugin_regFile[7][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][3]  ( .D(n4399), .CP(n7136), .Q(
        \RegFilePlugin_regFile[6][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][3]  ( .D(n4367), .CP(n7140), .Q(
        \RegFilePlugin_regFile[5][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][3]  ( .D(n4335), .CP(n7250), .Q(
        \RegFilePlugin_regFile[4][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][3]  ( .D(n4303), .CP(n7133), .Q(
        \RegFilePlugin_regFile[3][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][3]  ( .D(n4271), .CP(n7250), .Q(
        \RegFilePlugin_regFile[2][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][3]  ( .D(n4239), .CP(n7250), .Q(
        \RegFilePlugin_regFile[1][3] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][3]  ( .D(n4150), .CP(n7136), .Q(
        \RegFilePlugin_regFile[0][3] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[3]  ( .D(N851), .CP(n7134), .Q(
        _zz_RegFilePlugin_regFile_port0[3]) );
  dfnrq1 \decode_to_execute_RS1_reg[3]  ( .D(n4149), .CP(n7250), .Q(
        execute_RS1[3]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[3]  ( .D(N884), .CP(n7136), .Q(
        _zz_RegFilePlugin_regFile_port1[3]) );
  dfnrq1 \decode_to_execute_RS2_reg[3]  ( .D(n4148), .CP(n7134), .Q(
        execute_RS2[3]) );
  dfnrq1 \RegFilePlugin_regFile_reg[31][2]  ( .D(n5198), .CP(n7133), .Q(
        \RegFilePlugin_regFile[31][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[30][2]  ( .D(n5166), .CP(n7141), .Q(
        \RegFilePlugin_regFile[30][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[29][2]  ( .D(n5134), .CP(n7141), .Q(
        \RegFilePlugin_regFile[29][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[28][2]  ( .D(n5102), .CP(n7141), .Q(
        \RegFilePlugin_regFile[28][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[27][2]  ( .D(n5070), .CP(n7141), .Q(
        \RegFilePlugin_regFile[27][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[26][2]  ( .D(n5038), .CP(n7141), .Q(
        \RegFilePlugin_regFile[26][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[25][2]  ( .D(n5006), .CP(n7141), .Q(
        \RegFilePlugin_regFile[25][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[24][2]  ( .D(n4974), .CP(n7141), .Q(
        \RegFilePlugin_regFile[24][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[23][2]  ( .D(n4942), .CP(n7141), .Q(
        \RegFilePlugin_regFile[23][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[22][2]  ( .D(n4910), .CP(n7140), .Q(
        \RegFilePlugin_regFile[22][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[21][2]  ( .D(n4878), .CP(n7140), .Q(
        \RegFilePlugin_regFile[21][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[20][2]  ( .D(n4846), .CP(n7140), .Q(
        \RegFilePlugin_regFile[20][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[19][2]  ( .D(n4814), .CP(n7140), .Q(
        \RegFilePlugin_regFile[19][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[18][2]  ( .D(n4782), .CP(n7140), .Q(
        \RegFilePlugin_regFile[18][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[17][2]  ( .D(n4750), .CP(n7140), .Q(
        \RegFilePlugin_regFile[17][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[16][2]  ( .D(n4718), .CP(n7140), .Q(
        \RegFilePlugin_regFile[16][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[15][2]  ( .D(n4686), .CP(n7140), .Q(
        \RegFilePlugin_regFile[15][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[14][2]  ( .D(n4654), .CP(n7137), .Q(
        \RegFilePlugin_regFile[14][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[13][2]  ( .D(n4622), .CP(n7137), .Q(
        \RegFilePlugin_regFile[13][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[12][2]  ( .D(n4590), .CP(n7137), .Q(
        \RegFilePlugin_regFile[12][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[11][2]  ( .D(n4558), .CP(n7251), .Q(
        \RegFilePlugin_regFile[11][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[10][2]  ( .D(n4526), .CP(n7137), .Q(
        \RegFilePlugin_regFile[10][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[9][2]  ( .D(n4494), .CP(n7251), .Q(
        \RegFilePlugin_regFile[9][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[8][2]  ( .D(n4462), .CP(n7137), .Q(
        \RegFilePlugin_regFile[8][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[7][2]  ( .D(n4430), .CP(n7251), .Q(
        \RegFilePlugin_regFile[7][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[6][2]  ( .D(n4398), .CP(n7135), .Q(
        \RegFilePlugin_regFile[6][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[5][2]  ( .D(n4366), .CP(n7135), .Q(
        \RegFilePlugin_regFile[5][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[4][2]  ( .D(n4334), .CP(n7135), .Q(
        \RegFilePlugin_regFile[4][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[3][2]  ( .D(n4302), .CP(n7141), .Q(
        \RegFilePlugin_regFile[3][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[2][2]  ( .D(n4270), .CP(n7135), .Q(
        \RegFilePlugin_regFile[2][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[1][2]  ( .D(n4238), .CP(n7141), .Q(
        \RegFilePlugin_regFile[1][2] ) );
  dfnrq1 \RegFilePlugin_regFile_reg[0][2]  ( .D(n4147), .CP(n7135), .Q(
        \RegFilePlugin_regFile[0][2] ) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port0_reg[2]  ( .D(N852), .CP(n7141), .Q(
        _zz_RegFilePlugin_regFile_port0[2]) );
  dfnrq1 \decode_to_execute_RS1_reg[2]  ( .D(n4146), .CP(n7262), .Q(
        execute_RS1[2]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[2]  ( .D(N885), .CP(n7139), .Q(
        _zz_RegFilePlugin_regFile_port1[2]) );
  dfnrq1 \decode_to_execute_RS2_reg[2]  ( .D(n4145), .CP(n7262), .Q(
        execute_RS2[2]) );
  dfnrq1 \_zz_RegFilePlugin_regFile_port1_reg[1]  ( .D(N886), .CP(n7251), .Q(
        _zz_RegFilePlugin_regFile_port1[1]) );
  dfnrq1 \decode_to_execute_RS2_reg[1]  ( .D(n4142), .CP(n7262), .Q(
        execute_RS2[1]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[5]  ( .D(n6114), .CP(n7262), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[5]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[5]  ( 
        .D(n5240), .CP(n7262), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[5]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[5]  ( .D(
        n6180), .CP(n7141), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[5]) );
  dfnrq1 \CsrPlugin_mtval_reg[5]  ( .D(n6012), .CP(n7262), .Q(
        CsrPlugin_mtval[5]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[5]  ( .D(n6138), .CP(n7262), .Q(_zz_CsrPlugin_csrMapping_readDataInit[5]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[3]  ( .D(n4138), .CP(n7262), .Q(
        CsrPlugin_mtvec_base[3]) );
  dfnrq1 \decode_to_execute_PC_reg[5]  ( .D(n5239), .CP(n7262), .Q(
        execute_PC[5]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[5]  ( .D(n6067), .CP(n7137), .Q(
        debug_bus_rsp_data[5]) );
  dfnrq1 \memory_to_writeBack_PC_reg[3]  ( .D(n5232), .CP(n7251), .Q(
        writeBack_PC[3]) );
  dfnrq1 \CsrPlugin_mepc_reg[3]  ( .D(n4108), .CP(n7262), .Q(CsrPlugin_mepc[3]) );
  dfnrq1 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory_reg ( .D(N1783), .CP(n7262), .Q(CsrPlugin_exceptionPendings_2) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][2]  ( .D(n5325), .CP(n7251), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/banks_0_reg[0][1]  ( .D(n5324), .CP(n7251), 
        .Q(\IBusCachedPlugin_cache/banks_0[0][1] ) );
  dfnrq1 CsrPlugin_pipelineLiberator_pcValids_0_reg ( .D(n6131), .CP(n7138), 
        .Q(CsrPlugin_pipelineLiberator_pcValids_0) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_flushPending_reg  ( .D(n6081), 
        .CP(n7251), .Q(\IBusCachedPlugin_cache/lineLoader_flushPending ) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_flushCounter_reg[1]  ( .D(n6086), 
        .CP(n7138), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port[0] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_when_InstructionCache_l342_reg  ( .D(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port[0] ), .CP(n7250), .Q(
        \IBusCachedPlugin_cache/_zz_when_InstructionCache_l342 ) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_flushCounter_reg[0]  ( .D(n6087), 
        .CP(n7139), .Q(\IBusCachedPlugin_cache/lineLoader_flushCounter[0] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][0]  ( .D(n5888), .CP(n7251), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][27]  ( .D(n5887), .CP(
        n7251), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][26]  ( .D(n5886), .CP(
        n7250), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][25]  ( .D(n5885), .CP(
        n7141), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][24]  ( .D(n5884), .CP(
        n7134), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][23]  ( .D(n5883), .CP(
        n7251), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][22]  ( .D(n5882), .CP(
        n7250), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][21]  ( .D(n5881), .CP(
        n7251), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][20]  ( .D(n5880), .CP(
        n7133), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][19]  ( .D(n5879), .CP(
        n7251), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][18]  ( .D(n5878), .CP(
        n7251), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][17]  ( .D(n5877), .CP(
        n7135), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][16]  ( .D(n5876), .CP(
        n7137), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][15]  ( .D(n5875), .CP(
        n7140), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][14]  ( .D(n5874), .CP(
        n7141), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][13]  ( .D(n5873), .CP(
        n7135), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][12]  ( .D(n5872), .CP(
        n7137), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][11]  ( .D(n5871), .CP(
        n7139), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][10]  ( .D(n5870), .CP(
        n7139), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][9]  ( .D(n5869), .CP(n7139), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][8]  ( .D(n5868), .CP(n7139), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][7]  ( .D(n5867), .CP(n7139), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][6]  ( .D(n5866), .CP(n7139), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][5]  ( .D(n5865), .CP(n7139), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][4]  ( .D(n5864), .CP(n7139), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][3]  ( .D(n5863), .CP(n7138), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[1][2]  ( .D(n5862), .CP(n7138), .Q(\IBusCachedPlugin_cache/ways_0_tags[1][2] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][0]  ( .D(n5861), .CP(n7138), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][0] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][27]  ( .D(n5860), .CP(
        n7138), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][27] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][26]  ( .D(n5859), .CP(
        n7138), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][26] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][25]  ( .D(n5858), .CP(
        n7138), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][25] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][24]  ( .D(n5857), .CP(
        n7138), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][24] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][23]  ( .D(n5856), .CP(
        n7138), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][23] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][22]  ( .D(n5855), .CP(
        n7137), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][22] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][21]  ( .D(n5854), .CP(
        n7137), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][21] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][20]  ( .D(n5853), .CP(
        n7137), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][20] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][19]  ( .D(n5852), .CP(
        n7137), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][19] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][18]  ( .D(n5851), .CP(
        n7137), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][18] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][17]  ( .D(n5850), .CP(
        n7137), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][17] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][16]  ( .D(n5849), .CP(
        n7137), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][16] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][15]  ( .D(n5848), .CP(
        n7137), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][15] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][14]  ( .D(n5847), .CP(
        n7141), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][14] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][13]  ( .D(n5846), .CP(
        n7134), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][13] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][12]  ( .D(n5845), .CP(
        n7138), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][12] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][11]  ( .D(n5844), .CP(
        n7262), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][11] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][10]  ( .D(n5843), .CP(
        n7250), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][10] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][9]  ( .D(n5842), .CP(n7140), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][9] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][8]  ( .D(n5841), .CP(n7139), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][8] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][7]  ( .D(n5840), .CP(n7133), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][7] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][6]  ( .D(n5839), .CP(n7136), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][6] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][5]  ( .D(n5838), .CP(n7136), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][5] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][4]  ( .D(n5837), .CP(n7136), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][4] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][3]  ( .D(n5836), .CP(n7136), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][3] ) );
  dfnrq1 \IBusCachedPlugin_cache/ways_0_tags_reg[0][2]  ( .D(n5835), .CP(n7136), .Q(\IBusCachedPlugin_cache/ways_0_tags[0][2] ) );
  dfnrq1 DebugPlugin_haltedByBreak_reg ( .D(n6077), .CP(n7136), .Q(
        DebugPlugin_haltedByBreak) );
  dfnrq1 CsrPlugin_pipelineLiberator_pcValids_1_reg ( .D(n6132), .CP(n7136), 
        .Q(CsrPlugin_pipelineLiberator_pcValids_1) );
  dfnrq1 CsrPlugin_pipelineLiberator_pcValids_2_reg ( .D(n6133), .CP(n7136), 
        .Q(CsrPlugin_pipelineLiberator_pcValids_2) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[1]  ( .D(
        n6244), .CP(n7250), .Q(_zz_decode_LEGAL_INSTRUCTION_1[1]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[1]  ( .D(n5916), .CP(n7138), .Q(
        execute_INSTRUCTION[1]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[1]  ( .D(
        n6176), .CP(n7134), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[1]) );
  dfnrq1 \CsrPlugin_mtval_reg[1]  ( .D(n6008), .CP(n7134), .Q(
        CsrPlugin_mtval[1]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[4]  ( .D(n6115), .CP(n7133), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[4]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[4]  ( 
        .D(n5237), .CP(n7140), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[4]) );
  dfnrq1 \CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr_reg[4]  ( .D(
        n6179), .CP(n7139), .Q(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[4]) );
  dfnrq1 \CsrPlugin_mtval_reg[4]  ( .D(n6011), .CP(n7135), .Q(
        CsrPlugin_mtval[4]) );
  dfnrq1 \decode_to_execute_PC_reg[4]  ( .D(n5236), .CP(n7141), .Q(
        execute_PC[4]) );
  dfnrq1 \memory_to_writeBack_PC_reg[4]  ( .D(n5235), .CP(n7138), .Q(
        writeBack_PC[4]) );
  dfnrq1 \CsrPlugin_mepc_reg[4]  ( .D(n4107), .CP(n7262), .Q(CsrPlugin_mepc[4]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[4]  ( .D(n6137), .CP(n7134), .Q(_zz_CsrPlugin_csrMapping_readDataInit[4]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[2]  ( .D(n4139), .CP(n7133), .Q(
        CsrPlugin_mtvec_base[2]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[4]  ( .D(n6068), .CP(n7140), .Q(
        DebugPlugin_busReadDataReg[4]) );
  dfnrq1 \CsrPlugin_mcause_exceptionCode_reg[0]  ( .D(n4077), .CP(n7139), .Q(
        CsrPlugin_mcause_exceptionCode[0]) );
  dfnrq1 \CsrPlugin_mcause_exceptionCode_reg[1]  ( .D(n4076), .CP(n7135), .Q(
        CsrPlugin_mcause_exceptionCode[1]) );
  dfnrq1 \CsrPlugin_mepc_reg[1]  ( .D(n4110), .CP(n7136), .Q(CsrPlugin_mepc[1]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[1]  ( .D(n6134), .CP(n7139), .Q(_zz_CsrPlugin_csrMapping_readDataInit[1]) );
  dfnrq1 \CsrPlugin_mcause_exceptionCode_reg[2]  ( .D(n4075), .CP(n7140), .Q(
        CsrPlugin_mcause_exceptionCode[2]) );
  dfnrq1 \_zz_CsrPlugin_csrMapping_readDataInit_reg[2]  ( .D(n6135), .CP(n7133), .Q(_zz_CsrPlugin_csrMapping_readDataInit[2]) );
  dfnrq1 \CsrPlugin_mtvec_base_reg[0]  ( .D(n4141), .CP(n7134), .Q(
        CsrPlugin_mtvec_base[0]) );
  dfnrq1 IBusCachedPlugin_fetchPc_inc_reg ( .D(n6118), .CP(n7138), .Q(
        \_zz_IBusCachedPlugin_fetchPc_pc_1[2] ) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[0]  ( .D(n5977), .CP(n7251), .Q(
        execute_INSTRUCTION[0]) );
  dfnrq1 \IBusCachedPlugin_fetchPc_pcReg_reg[2]  ( .D(n6117), .CP(n7139), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[2]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[2]  ( .D(n6070), .CP(n7135), .Q(
        DebugPlugin_busReadDataReg[2]) );
  dfnrq1 \_zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload_reg[12]  ( 
        .D(n5261), .CP(n7135), .Q(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[12]) );
  dfnrq1 \decode_to_execute_PC_reg[12]  ( .D(n5260), .CP(n7135), .Q(
        execute_PC[12]) );
  dfnrq1 \memory_to_writeBack_PC_reg[12]  ( .D(n5259), .CP(n7135), .Q(
        writeBack_PC[12]) );
  dfnrq1 \CsrPlugin_mepc_reg[12]  ( .D(n4099), .CP(n7135), .Q(
        CsrPlugin_mepc[12]) );
  dfnrq1 \DebugPlugin_busReadDataReg_reg[12]  ( .D(n6060), .CP(n7135), .Q(
        debug_bus_rsp_data[12]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[31]  ( .D(n4067), .CP(
        n7135), .Q(\IBusCachedPlugin_cache/n2 ) );
  dfnrq1 execute_to_memory_BRANCH_DO_reg ( .D(n4066), .CP(n7135), .Q(
        memory_BRANCH_DO) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_hit_valid_reg  ( .D(n4065), .CP(
        n7134), .Q(\IBusCachedPlugin_cache/decodeStage_hit_valid ) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[12]  ( 
        .D(n4064), .CP(n7134), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[12]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[30]  ( 
        .D(n4063), .CP(n7134), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[30]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[31]  ( 
        .D(n4062), .CP(n7134), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[31]) );
  dfnrq1 \execute_to_memory_PC_reg[2]  ( .D(n4060), .CP(n7134), .Q(
        memory_PC[2]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[0]  ( .D(n4059), .CP(
        n7134), .Q(\IBusCachedPlugin_cache/n23 ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[2]  ( .D(n4058), .CP(
        n7134), .Q(\IBusCachedPlugin_cache/n21 ) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[31]  ( .D(n4057), .CP(n7134), .Q(
        memory_BRANCH_CALC[31]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[30]  ( .D(n4056), .CP(n7133), .Q(
        memory_BRANCH_CALC[30]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[29]  ( .D(n4055), .CP(n7136), .Q(
        memory_BRANCH_CALC[29]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[28]  ( .D(n4054), .CP(n7140), .Q(
        memory_BRANCH_CALC[28]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[27]  ( .D(n4053), .CP(n7136), .Q(
        memory_BRANCH_CALC[27]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[26]  ( .D(n4052), .CP(n7139), .Q(
        memory_BRANCH_CALC[26]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[25]  ( .D(n4051), .CP(n7136), .Q(
        memory_BRANCH_CALC[25]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[24]  ( .D(n4050), .CP(n7135), .Q(
        memory_BRANCH_CALC[24]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[23]  ( .D(n4049), .CP(n7136), .Q(
        memory_BRANCH_CALC[23]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[22]  ( .D(n4048), .CP(n7133), .Q(
        memory_BRANCH_CALC[22]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[21]  ( .D(n4047), .CP(n7133), .Q(
        memory_BRANCH_CALC[21]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[20]  ( .D(n4046), .CP(n7133), .Q(
        memory_BRANCH_CALC[20]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[19]  ( .D(n4045), .CP(n7133), .Q(
        memory_BRANCH_CALC[19]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[18]  ( .D(n4044), .CP(n7133), .Q(
        memory_BRANCH_CALC[18]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[17]  ( .D(n4043), .CP(n7133), .Q(
        memory_BRANCH_CALC[17]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[16]  ( .D(n4042), .CP(n7133), .Q(
        memory_BRANCH_CALC[16]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[15]  ( .D(n4041), .CP(n7133), .Q(
        memory_BRANCH_CALC[15]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[14]  ( .D(n4040), .CP(n7128), .Q(
        memory_BRANCH_CALC[14]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[13]  ( .D(n4039), .CP(n7127), .Q(
        memory_BRANCH_CALC[13]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[12]  ( .D(n4038), .CP(n7263), .Q(
        memory_BRANCH_CALC[12]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[11]  ( .D(n4037), .CP(n7125), .Q(
        memory_BRANCH_CALC[11]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[10]  ( .D(n4036), .CP(n7124), .Q(
        memory_BRANCH_CALC[10]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[9]  ( .D(n4035), .CP(n7128), .Q(
        memory_BRANCH_CALC[9]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[8]  ( .D(n4034), .CP(n7126), .Q(
        memory_BRANCH_CALC[8]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[7]  ( .D(n4033), .CP(n7129), .Q(
        memory_BRANCH_CALC[7]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[6]  ( .D(n4032), .CP(n7132), .Q(
        memory_BRANCH_CALC[6]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[5]  ( .D(n4031), .CP(n7132), .Q(
        memory_BRANCH_CALC[5]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[4]  ( .D(n4030), .CP(n7132), .Q(
        memory_BRANCH_CALC[4]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[3]  ( .D(n4029), .CP(n7132), .Q(
        memory_BRANCH_CALC[3]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[2]  ( .D(n4028), .CP(n7132), .Q(
        memory_BRANCH_CALC[2]) );
  dfnrq1 \execute_to_memory_BRANCH_CALC_reg[1]  ( .D(n4027), .CP(n7132), .Q(
        memory_BRANCH_CALC[1]) );
  dfnrq1 \execute_to_memory_PC_reg[31]  ( .D(n4025), .CP(n7132), .Q(
        memory_PC[31]) );
  dfnrq1 \execute_to_memory_PC_reg[30]  ( .D(n4024), .CP(n7132), .Q(
        memory_PC[30]) );
  dfnrq1 \execute_to_memory_PC_reg[3]  ( .D(n4023), .CP(n7130), .Q(
        memory_PC[3]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[3]  ( .D(n4021), .CP(
        n7132), .Q(\IBusCachedPlugin_cache/n20 ) );
  dfnrq1 execute_to_memory_MEMORY_ENABLE_reg ( .D(n4020), .CP(n7127), .Q(
        memory_MEMORY_ENABLE) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[30]  ( .D(n4019), .CP(
        n7129), .Q(\IBusCachedPlugin_cache/n3 ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[29]  ( .D(n4018), .CP(
        n7263), .Q(\IBusCachedPlugin_cache/n4 ) );
  dfnrq1 \execute_to_memory_INSTRUCTION_reg[29]  ( .D(n4017), .CP(clk), .Q(
        memory_INSTRUCTION_29) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[28]  ( .D(n4016), .CP(
        n7128), .Q(\IBusCachedPlugin_cache/n5 ) );
  dfnrq1 \execute_to_memory_INSTRUCTION_reg[28]  ( .D(n4015), .CP(n7125), .Q(
        memory_INSTRUCTION_28) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[27]  ( .D(n4014), .CP(
        n7263), .Q(\IBusCachedPlugin_cache/n6 ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[26]  ( .D(n4013), .CP(
        n7131), .Q(\IBusCachedPlugin_cache/n7 ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[25]  ( .D(n4012), .CP(
        n7263), .Q(\IBusCachedPlugin_cache/n8 ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[24]  ( .D(n4011), .CP(
        n7126), .Q(IBusCachedPlugin_cache_io_cpu_fetch_data[24]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[23]  ( .D(n4010), .CP(
        n7263), .Q(IBusCachedPlugin_cache_io_cpu_fetch_data[23]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[22]  ( .D(n4009), .CP(
        n7130), .Q(IBusCachedPlugin_cache_io_cpu_fetch_data[22]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[21]  ( .D(n4008), .CP(
        n7263), .Q(IBusCachedPlugin_cache_io_cpu_fetch_data[21]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[20]  ( .D(n4007), .CP(
        n7132), .Q(IBusCachedPlugin_cache_io_cpu_fetch_data[20]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[19]  ( .D(n4006), .CP(
        n7132), .Q(IBusCachedPlugin_cache_io_cpu_fetch_data[19]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[18]  ( .D(n4005), .CP(
        n7129), .Q(IBusCachedPlugin_cache_io_cpu_fetch_data[18]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[17]  ( .D(n4004), .CP(
        n7130), .Q(IBusCachedPlugin_cache_io_cpu_fetch_data[17]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[16]  ( .D(n4003), .CP(
        n7131), .Q(IBusCachedPlugin_cache_io_cpu_fetch_data[16]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[15]  ( .D(n4002), .CP(
        n7126), .Q(IBusCachedPlugin_cache_io_cpu_fetch_data[15]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[14]  ( .D(n4001), .CP(
        n7130), .Q(\IBusCachedPlugin_cache/n9 ) );
  dfnrq1 \execute_to_memory_INSTRUCTION_reg[14]  ( .D(n4000), .CP(n7132), .Q(
        memory_INSTRUCTION[14]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[13]  ( .D(n3999), .CP(
        n7129), .Q(\IBusCachedPlugin_cache/n10 ) );
  dfnrq1 \dBus_cmd_rData_size_reg[1]  ( .D(n3998), .CP(n7131), .Q(
        dBus_cmd_halfPipe_payload_size[1]) );
  dfnrq1 \execute_to_memory_INSTRUCTION_reg[13]  ( .D(n3997), .CP(n7131), .Q(
        memory_INSTRUCTION[13]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[12]  ( .D(n3996), .CP(
        n7131), .Q(\IBusCachedPlugin_cache/n11 ) );
  dfnrq1 \execute_to_memory_INSTRUCTION_reg[12]  ( .D(n3995), .CP(n7131), .Q(
        memory_INSTRUCTION[12]) );
  dfnrq1 \dBus_cmd_rData_size_reg[0]  ( .D(n3994), .CP(n7131), .Q(
        dBus_cmd_halfPipe_payload_size[0]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[11]  ( .D(n3993), .CP(
        n7131), .Q(\IBusCachedPlugin_cache/n12 ) );
  dfnrq1 \execute_to_memory_INSTRUCTION_reg[11]  ( .D(n3992), .CP(n7131), .Q(
        memory_INSTRUCTION[11]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[10]  ( .D(n3991), .CP(
        n7131), .Q(\IBusCachedPlugin_cache/n13 ) );
  dfnrq1 \execute_to_memory_INSTRUCTION_reg[10]  ( .D(n3990), .CP(n7123), .Q(
        memory_INSTRUCTION[10]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[9]  ( .D(n3989), .CP(
        n7124), .Q(\IBusCachedPlugin_cache/n14 ) );
  dfnrq1 \execute_to_memory_INSTRUCTION_reg[9]  ( .D(n3988), .CP(n7123), .Q(
        memory_INSTRUCTION[9]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[8]  ( .D(n3987), .CP(
        n7124), .Q(\IBusCachedPlugin_cache/n15 ) );
  dfnrq1 \execute_to_memory_INSTRUCTION_reg[8]  ( .D(n3986), .CP(n7123), .Q(
        memory_INSTRUCTION[8]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[7]  ( .D(n3985), .CP(
        n7124), .Q(\IBusCachedPlugin_cache/n16 ) );
  dfnrq1 \execute_to_memory_INSTRUCTION_reg[7]  ( .D(n3984), .CP(n7123), .Q(
        memory_INSTRUCTION[7]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[6]  ( .D(n3983), .CP(
        n7124), .Q(\IBusCachedPlugin_cache/n17 ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[5]  ( .D(n3982), .CP(
        n7125), .Q(\IBusCachedPlugin_cache/n18 ) );
  dfnrq1 execute_to_memory_MEMORY_STORE_reg ( .D(n3981), .CP(n7263), .Q(
        memory_MEMORY_STORE) );
  dfnrq1 dBus_cmd_rData_wr_reg ( .D(n3980), .CP(n7132), .Q(dBusWishbone_WE) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[4]  ( .D(n3979), .CP(
        n7127), .Q(\IBusCachedPlugin_cache/n19 ) );
  dfnrq1 \execute_to_memory_ENV_CTRL_reg[0]  ( .D(n3978), .CP(n7126), .Q(
        memory_ENV_CTRL[0]) );
  dfnrq1 \execute_to_memory_ENV_CTRL_reg[1]  ( .D(n3977), .CP(n7129), .Q(
        memory_ENV_CTRL[1]) );
  dfnrq1 execute_to_memory_REGFILE_WRITE_VALID_reg ( .D(n3976), .CP(n7130), 
        .Q(memory_REGFILE_WRITE_VALID) );
  dfnrq1 \execute_to_memory_MEMORY_ADDRESS_LOW_reg[0]  ( .D(n3975), .CP(n7124), 
        .Q(memory_MEMORY_ADDRESS_LOW[0]) );
  dfnrq1 \execute_to_memory_MEMORY_ADDRESS_LOW_reg[1]  ( .D(n3974), .CP(n7124), 
        .Q(memory_MEMORY_ADDRESS_LOW[1]) );
  dfnrq1 \dBus_cmd_rData_data_reg[0]  ( .D(n3973), .CP(n7125), .Q(
        dBusWishbone_DAT_MOSI[0]) );
  dfnrq1 \dBus_cmd_rData_address_reg[31]  ( .D(n3972), .CP(n7130), .Q(
        dBusWishbone_ADR[29]) );
  dfnrq1 \dBus_cmd_rData_address_reg[30]  ( .D(n3971), .CP(n7125), .Q(
        dBusWishbone_ADR[28]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[29]  ( 
        .D(n3970), .CP(n7128), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[29]) );
  dfnrq1 \execute_to_memory_PC_reg[29]  ( .D(n3969), .CP(n7130), .Q(
        memory_PC[29]) );
  dfnrq1 \dBus_cmd_rData_address_reg[29]  ( .D(n3968), .CP(n7125), .Q(
        dBusWishbone_ADR[27]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[28]  ( 
        .D(n3967), .CP(n7132), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[28]) );
  dfnrq1 \execute_to_memory_PC_reg[28]  ( .D(n3966), .CP(n7130), .Q(
        memory_PC[28]) );
  dfnrq1 \dBus_cmd_rData_address_reg[28]  ( .D(n3965), .CP(n7130), .Q(
        dBusWishbone_ADR[26]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[27]  ( 
        .D(n3964), .CP(n7130), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[27]) );
  dfnrq1 \execute_to_memory_PC_reg[27]  ( .D(n3963), .CP(n7130), .Q(
        memory_PC[27]) );
  dfnrq1 \dBus_cmd_rData_address_reg[27]  ( .D(n3962), .CP(n7130), .Q(
        dBusWishbone_ADR[25]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[26]  ( 
        .D(n3961), .CP(n7130), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[26]) );
  dfnrq1 \execute_to_memory_PC_reg[26]  ( .D(n3960), .CP(n7130), .Q(
        memory_PC[26]) );
  dfnrq1 \dBus_cmd_rData_address_reg[26]  ( .D(n3959), .CP(n7130), .Q(
        dBusWishbone_ADR[24]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[25]  ( 
        .D(n3958), .CP(n7129), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[25]) );
  dfnrq1 \execute_to_memory_PC_reg[25]  ( .D(n3957), .CP(n7129), .Q(
        memory_PC[25]) );
  dfnrq1 \dBus_cmd_rData_address_reg[25]  ( .D(n3956), .CP(n7129), .Q(
        dBusWishbone_ADR[23]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[24]  ( 
        .D(n3955), .CP(n7129), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[24]) );
  dfnrq1 \execute_to_memory_PC_reg[24]  ( .D(n3954), .CP(n7129), .Q(
        memory_PC[24]) );
  dfnrq1 \dBus_cmd_rData_address_reg[24]  ( .D(n3953), .CP(n7129), .Q(
        dBusWishbone_ADR[22]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[23]  ( 
        .D(n3952), .CP(n7129), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[23]) );
  dfnrq1 \execute_to_memory_PC_reg[23]  ( .D(n3951), .CP(n7129), .Q(
        memory_PC[23]) );
  dfnrq1 \dBus_cmd_rData_address_reg[23]  ( .D(n3950), .CP(n7123), .Q(
        dBusWishbone_ADR[21]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[22]  ( 
        .D(n3949), .CP(n7123), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[22]) );
  dfnrq1 \execute_to_memory_PC_reg[22]  ( .D(n3948), .CP(n7123), .Q(
        memory_PC[22]) );
  dfnrq1 \dBus_cmd_rData_address_reg[22]  ( .D(n3947), .CP(n7123), .Q(
        dBusWishbone_ADR[20]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[21]  ( 
        .D(n3946), .CP(n7123), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[21]) );
  dfnrq1 \execute_to_memory_PC_reg[21]  ( .D(n3945), .CP(n7123), .Q(
        memory_PC[21]) );
  dfnrq1 \dBus_cmd_rData_address_reg[21]  ( .D(n3944), .CP(n7123), .Q(
        dBusWishbone_ADR[19]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[20]  ( 
        .D(n3943), .CP(n7123), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[20]) );
  dfnrq1 \execute_to_memory_PC_reg[20]  ( .D(n3942), .CP(n7126), .Q(
        memory_PC[20]) );
  dfnrq1 \dBus_cmd_rData_address_reg[20]  ( .D(n3941), .CP(n7131), .Q(
        dBusWishbone_ADR[18]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[19]  ( 
        .D(n3940), .CP(n7131), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[19]) );
  dfnrq1 \execute_to_memory_PC_reg[19]  ( .D(n3939), .CP(n7132), .Q(
        memory_PC[19]) );
  dfnrq1 \dBus_cmd_rData_address_reg[19]  ( .D(n3938), .CP(n7263), .Q(
        dBusWishbone_ADR[17]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[18]  ( 
        .D(n3937), .CP(n7263), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[18]) );
  dfnrq1 \execute_to_memory_PC_reg[18]  ( .D(n3936), .CP(n7129), .Q(
        memory_PC[18]) );
  dfnrq1 \dBus_cmd_rData_address_reg[18]  ( .D(n3935), .CP(n7125), .Q(
        dBusWishbone_ADR[16]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[17]  ( 
        .D(n3934), .CP(n7123), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[17]) );
  dfnrq1 \execute_to_memory_PC_reg[17]  ( .D(n3933), .CP(n7123), .Q(
        memory_PC[17]) );
  dfnrq1 \dBus_cmd_rData_address_reg[17]  ( .D(n3932), .CP(n7128), .Q(
        dBusWishbone_ADR[15]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[16]  ( 
        .D(n3931), .CP(n7127), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[16]) );
  dfnrq1 \execute_to_memory_PC_reg[16]  ( .D(n3930), .CP(n7132), .Q(
        memory_PC[16]) );
  dfnrq1 \dBus_cmd_rData_address_reg[16]  ( .D(n3929), .CP(n7124), .Q(
        dBusWishbone_ADR[14]) );
  dfnrq1 \dBus_cmd_rData_data_reg[16]  ( .D(n3928), .CP(n7127), .Q(
        dBusWishbone_DAT_MOSI[16]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[15]  ( 
        .D(n3927), .CP(n7123), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[15]) );
  dfnrq1 \execute_to_memory_PC_reg[15]  ( .D(n3926), .CP(n7128), .Q(
        memory_PC[15]) );
  dfnrq1 \dBus_cmd_rData_address_reg[15]  ( .D(n3925), .CP(n7128), .Q(
        dBusWishbone_ADR[13]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[14]  ( 
        .D(n3924), .CP(n7128), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[14]) );
  dfnrq1 \execute_to_memory_PC_reg[14]  ( .D(n3923), .CP(n7128), .Q(
        memory_PC[14]) );
  dfnrq1 \dBus_cmd_rData_address_reg[14]  ( .D(n3922), .CP(n7128), .Q(
        dBusWishbone_ADR[12]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[13]  ( 
        .D(n3921), .CP(n7128), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[13]) );
  dfnrq1 \execute_to_memory_PC_reg[13]  ( .D(n3920), .CP(n7128), .Q(
        memory_PC[13]) );
  dfnrq1 \dBus_cmd_rData_address_reg[13]  ( .D(n3919), .CP(n7128), .Q(
        dBusWishbone_ADR[11]) );
  dfnrq1 \dBus_cmd_rData_address_reg[12]  ( .D(n3918), .CP(n7125), .Q(
        dBusWishbone_ADR[10]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[11]  ( 
        .D(n3917), .CP(n7131), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[11]) );
  dfnrq1 \execute_to_memory_PC_reg[11]  ( .D(n3916), .CP(n7126), .Q(
        memory_PC[11]) );
  dfnrq1 \dBus_cmd_rData_address_reg[11]  ( .D(n3915), .CP(n7129), .Q(
        dBusWishbone_ADR[9]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[10]  ( 
        .D(n3914), .CP(n7263), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[10]) );
  dfnrq1 \execute_to_memory_PC_reg[10]  ( .D(n3913), .CP(n7131), .Q(
        memory_PC[10]) );
  dfnrq1 \dBus_cmd_rData_address_reg[10]  ( .D(n3912), .CP(n7263), .Q(
        dBusWishbone_ADR[8]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[9]  ( 
        .D(n3911), .CP(n7131), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[9]) );
  dfnrq1 \execute_to_memory_PC_reg[9]  ( .D(n3910), .CP(n7127), .Q(
        memory_PC[9]) );
  dfnrq1 \dBus_cmd_rData_address_reg[9]  ( .D(n3909), .CP(n7127), .Q(
        dBusWishbone_ADR[7]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[8]  ( 
        .D(n3908), .CP(n7127), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[8]) );
  dfnrq1 \execute_to_memory_PC_reg[8]  ( .D(n3907), .CP(n7127), .Q(
        memory_PC[8]) );
  dfnrq1 \dBus_cmd_rData_address_reg[8]  ( .D(n3906), .CP(n7127), .Q(
        dBusWishbone_ADR[6]) );
  dfnrq1 \dBus_cmd_rData_data_reg[8]  ( .D(n3905), .CP(n7127), .Q(
        dBusWishbone_DAT_MOSI[8]) );
  dfnrq1 \dBus_cmd_rData_data_reg[24]  ( .D(n3904), .CP(n7127), .Q(
        dBusWishbone_DAT_MOSI[24]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[7]  ( 
        .D(n3903), .CP(n7127), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[7]) );
  dfnrq1 \execute_to_memory_PC_reg[7]  ( .D(n3902), .CP(n7126), .Q(
        memory_PC[7]) );
  dfnrq1 \dBus_cmd_rData_address_reg[7]  ( .D(n3901), .CP(n7126), .Q(
        dBusWishbone_ADR[5]) );
  dfnrq1 \dBus_cmd_rData_data_reg[7]  ( .D(n3900), .CP(n7126), .Q(
        dBusWishbone_DAT_MOSI[7]) );
  dfnrq1 \dBus_cmd_rData_data_reg[15]  ( .D(n3899), .CP(n7126), .Q(
        dBusWishbone_DAT_MOSI[15]) );
  dfnrq1 \dBus_cmd_rData_data_reg[23]  ( .D(n3898), .CP(n7126), .Q(
        dBusWishbone_DAT_MOSI[23]) );
  dfnrq1 \dBus_cmd_rData_data_reg[31]  ( .D(n3897), .CP(n7126), .Q(
        dBusWishbone_DAT_MOSI[31]) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[6]  ( 
        .D(n3896), .CP(n7126), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[6]) );
  dfnrq1 \execute_to_memory_PC_reg[6]  ( .D(n3895), .CP(n7126), .Q(
        memory_PC[6]) );
  dfnrq1 \dBus_cmd_rData_address_reg[6]  ( .D(n3894), .CP(n7263), .Q(
        dBusWishbone_ADR[4]) );
  dfnrq1 \dBus_cmd_rData_data_reg[6]  ( .D(n3893), .CP(n7129), .Q(
        dBusWishbone_DAT_MOSI[6]) );
  dfnrq1 \dBus_cmd_rData_data_reg[14]  ( .D(n3892), .CP(n7130), .Q(
        dBusWishbone_DAT_MOSI[14]) );
  dfnrq1 \dBus_cmd_rData_data_reg[22]  ( .D(n3891), .CP(n7127), .Q(
        dBusWishbone_DAT_MOSI[22]) );
  dfnrq1 \dBus_cmd_rData_data_reg[30]  ( .D(n3890), .CP(n7126), .Q(
        dBusWishbone_DAT_MOSI[30]) );
  dfnrq1 \dBus_cmd_rData_address_reg[5]  ( .D(n3889), .CP(n7126), .Q(
        dBusWishbone_ADR[3]) );
  dfnrq1 \dBus_cmd_rData_data_reg[5]  ( .D(n3888), .CP(n7263), .Q(
        dBusWishbone_DAT_MOSI[5]) );
  dfnrq1 \dBus_cmd_rData_data_reg[13]  ( .D(n3887), .CP(n7131), .Q(
        dBusWishbone_DAT_MOSI[13]) );
  dfnrq1 \dBus_cmd_rData_data_reg[21]  ( .D(n3886), .CP(n7125), .Q(
        dBusWishbone_DAT_MOSI[21]) );
  dfnrq1 \dBus_cmd_rData_data_reg[29]  ( .D(n3885), .CP(n7125), .Q(
        dBusWishbone_DAT_MOSI[29]) );
  dfnrq1 \dBus_cmd_rData_address_reg[4]  ( .D(n3884), .CP(n7125), .Q(
        dBusWishbone_ADR[2]) );
  dfnrq1 \dBus_cmd_rData_data_reg[4]  ( .D(n3883), .CP(n7125), .Q(
        dBusWishbone_DAT_MOSI[4]) );
  dfnrq1 \dBus_cmd_rData_data_reg[12]  ( .D(n3882), .CP(n7125), .Q(
        dBusWishbone_DAT_MOSI[12]) );
  dfnrq1 \dBus_cmd_rData_data_reg[20]  ( .D(n3881), .CP(n7125), .Q(
        dBusWishbone_DAT_MOSI[20]) );
  dfnrq1 \dBus_cmd_rData_data_reg[28]  ( .D(n3880), .CP(n7125), .Q(
        dBusWishbone_DAT_MOSI[28]) );
  dfnrq1 \dBus_cmd_rData_address_reg[3]  ( .D(n3879), .CP(n7125), .Q(
        dBusWishbone_ADR[1]) );
  dfnrq1 \dBus_cmd_rData_data_reg[3]  ( .D(n3878), .CP(n7129), .Q(
        dBusWishbone_DAT_MOSI[3]) );
  dfnrq1 \dBus_cmd_rData_data_reg[11]  ( .D(n3877), .CP(n7125), .Q(
        dBusWishbone_DAT_MOSI[11]) );
  dfnrq1 \dBus_cmd_rData_data_reg[19]  ( .D(n3876), .CP(n7131), .Q(
        dBusWishbone_DAT_MOSI[19]) );
  dfnrq1 \dBus_cmd_rData_data_reg[27]  ( .D(n3875), .CP(n7126), .Q(
        dBusWishbone_DAT_MOSI[27]) );
  dfnrq1 \dBus_cmd_rData_address_reg[2]  ( .D(n3874), .CP(n7130), .Q(
        dBusWishbone_ADR[0]) );
  dfnrq1 \dBus_cmd_rData_data_reg[2]  ( .D(n3873), .CP(n7132), .Q(
        dBusWishbone_DAT_MOSI[2]) );
  dfnrq1 \dBus_cmd_rData_data_reg[10]  ( .D(n3872), .CP(n7129), .Q(
        dBusWishbone_DAT_MOSI[10]) );
  dfnrq1 \dBus_cmd_rData_data_reg[18]  ( .D(n3871), .CP(n7263), .Q(
        dBusWishbone_DAT_MOSI[18]) );
  dfnrq1 \dBus_cmd_rData_data_reg[26]  ( .D(n3870), .CP(n7263), .Q(
        dBusWishbone_DAT_MOSI[26]) );
  dfnrq1 \dBus_cmd_rData_address_reg[1]  ( .D(n3869), .CP(n7131), .Q(
        dBus_cmd_halfPipe_payload_address[1]) );
  dfnrq1 \dBus_cmd_rData_data_reg[1]  ( .D(n3868), .CP(n7126), .Q(
        dBusWishbone_DAT_MOSI[1]) );
  dfnrq1 \dBus_cmd_rData_data_reg[9]  ( .D(n3867), .CP(n7130), .Q(
        dBusWishbone_DAT_MOSI[9]) );
  dfnrq1 \dBus_cmd_rData_data_reg[17]  ( .D(n3866), .CP(n7132), .Q(
        dBusWishbone_DAT_MOSI[17]) );
  dfnrq1 \dBus_cmd_rData_data_reg[25]  ( .D(n3865), .CP(n7127), .Q(
        dBusWishbone_DAT_MOSI[25]) );
  dfnrq1 \dBus_cmd_rData_address_reg[0]  ( .D(n3864), .CP(n7263), .Q(
        dBus_cmd_halfPipe_payload_address[0]) );
  dfnrq1 execute_to_memory_ALIGNEMENT_FAULT_reg ( .D(n3863), .CP(n7129), .Q(
        memory_ALIGNEMENT_FAULT) );
  dfnrq1 \IBusCachedPlugin_cache/decodeStage_mmuRsp_physicalAddress_reg[5]  ( 
        .D(n3862), .CP(n7128), .Q(
        IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[5]) );
  dfnrq1 \execute_to_memory_PC_reg[5]  ( .D(n3861), .CP(n7127), .Q(
        memory_PC[5]) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[0]  ( .D(n3860), 
        .CP(n7128), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[0] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[27]  ( .D(n3859), 
        .CP(n7127), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[27] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[26]  ( .D(n3858), 
        .CP(n7128), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[26] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[25]  ( .D(n3857), 
        .CP(n7127), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[25] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[24]  ( .D(n3856), 
        .CP(n7128), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[24] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[23]  ( .D(n3855), 
        .CP(n7127), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[23] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[22]  ( .D(n3854), 
        .CP(n7124), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[22] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[21]  ( .D(n3853), 
        .CP(n7124), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[21] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[20]  ( .D(n3852), 
        .CP(n7124), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[20] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[19]  ( .D(n3851), 
        .CP(n7124), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[19] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[18]  ( .D(n3850), 
        .CP(n7124), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[18] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[17]  ( .D(n3849), 
        .CP(n7124), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[17] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[16]  ( .D(n3848), 
        .CP(n7124), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[16] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[15]  ( .D(n3847), 
        .CP(n7124), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[15] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[14]  ( .D(n3846), 
        .CP(n7123), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[14] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[13]  ( .D(n3845), 
        .CP(n7123), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[13] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[12]  ( .D(n3844), 
        .CP(n7123), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[12] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[11]  ( .D(n3843), 
        .CP(n7123), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[11] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[10]  ( .D(n3842), 
        .CP(n7123), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[10] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[9]  ( .D(n3841), 
        .CP(n7123), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[9] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[8]  ( .D(n3840), 
        .CP(n7123), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[8] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[7]  ( .D(n3839), 
        .CP(n7123), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[7] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[6]  ( .D(n3838), 
        .CP(n7263), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[6] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[5]  ( .D(n3837), 
        .CP(n7132), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[5] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[4]  ( .D(n3836), 
        .CP(n7131), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[4] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[3]  ( .D(n3835), 
        .CP(n7126), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[3] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_ways_0_tags_port1_reg[2]  ( .D(n3834), 
        .CP(n7125), .Q(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[2] ) );
  dfnrq1 \IBusCachedPlugin_cache/_zz_banks_0_port1_reg[1]  ( .D(n3833), .CP(
        n7130), .Q(\IBusCachedPlugin_cache/n22 ) );
  dfnrq1 \execute_to_memory_PC_reg[4]  ( .D(n3832), .CP(n7124), .Q(
        memory_PC[4]) );
  dfnrq1 \execute_to_memory_PC_reg[12]  ( .D(n3831), .CP(n7123), .Q(
        memory_PC[12]) );
  dfnrq1 \decode_to_execute_INSTRUCTION_reg[31]  ( .D(n5976), .CP(n7228), .Q(
        _zz__zz_execute_SRC2_3[11]) );
  dfnrq1 dBus_cmd_rValid_reg ( .D(n6175), .CP(n7230), .Q(n7265) );
  dfnrq1 \IBusCachedPlugin_cache/lineLoader_wordIndex_reg[2]  ( .D(n6083), 
        .CP(n7226), .Q(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[2] )
         );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[28]  ( .D(
        n6217), .CP(n7204), .Q(_zz_decode_LEGAL_INSTRUCTION_13[28]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[20]  ( .D(
        n6225), .CP(n7198), .Q(\_zz__zz_decode_ENV_CTRL_2_1[20] ) );
  dfnrq1 execute_CsrPlugin_csr_833_reg ( .D(n6003), .CP(n7198), .Q(
        execute_CsrPlugin_csr_833) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[14]  ( .D(
        n6231), .CP(n7237), .Q(\_zz_decode_LEGAL_INSTRUCTION_7[14] ) );
  dfnrq1 \memory_to_writeBack_INSTRUCTION_reg[9]  ( .D(memory_INSTRUCTION[9]), 
        .CP(n7237), .Q(_zz_lastStageRegFileWrite_payload_address[9]) );
  dfnrq1 \memory_to_writeBack_INSTRUCTION_reg[8]  ( .D(memory_INSTRUCTION[8]), 
        .CP(n7202), .Q(_zz_lastStageRegFileWrite_payload_address[8]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[6]  ( .D(
        n6239), .CP(n7201), .Q(_zz_decode_LEGAL_INSTRUCTION_1[6]) );
  dfnrq1 \IBusCachedPlugin_cache/io_cpu_fetch_data_regNextWhen_reg[4]  ( .D(
        n6241), .CP(n7201), .Q(_zz_decode_LEGAL_INSTRUCTION_1[4]) );
  dfnrb1 _zz_when_DebugPlugin_l244_reg ( .D(debug_bus_cmd_payload_address[2]), 
        .CP(n7229), .Q(_zz_when_DebugPlugin_l244), .QN(n7264) );
  inv0d1 U4 ( .I(n3250), .ZN(n3230) );
  aoi21d1 U5 ( .B1(debug_bus_cmd_payload_data[25]), .B2(n2429), .A(debugReset), 
        .ZN(n2433) );
  buffd1 U6 ( .I(n416), .Z(n531) );
  nr02d1 U7 ( .A1(n7007), .A2(n2094), .ZN(n2095) );
  inv0d1 U8 ( .I(iBus_rsp_payload_data[27]), .ZN(n3176) );
  inv0d1 U9 ( .I(iBus_rsp_payload_data[28]), .ZN(n3175) );
  inv0d1 U10 ( .I(iBus_rsp_payload_data[30]), .ZN(n3173) );
  inv0d1 U11 ( .I(iBus_rsp_payload_data[26]), .ZN(n3177) );
  inv0d1 U12 ( .I(n2086), .ZN(n2094) );
  inv0d1 U13 ( .I(iBus_rsp_payload_data[29]), .ZN(n3174) );
  inv0d1 U14 ( .I(iBus_rsp_payload_data[24]), .ZN(n3179) );
  inv0d1 U15 ( .I(n2749), .ZN(n3020) );
  inv0d1 U16 ( .I(n2356), .ZN(n6936) );
  inv0d4 U17 ( .I(n2135), .ZN(n2198) );
  nd02d2 U18 ( .A1(n313), .A2(n3679), .ZN(n314) );
  inv0d1 U19 ( .I(n3003), .ZN(n2932) );
  aoi22d1 U20 ( .A1(n2615), .A2(memory_INSTRUCTION[9]), .B1(n2614), .B2(
        memory_INSTRUCTION[10]), .ZN(n224) );
  nd02d2 U21 ( .A1(n6343), .A2(n308), .ZN(n305) );
  nr02d1 U22 ( .A1(n2996), .A2(n3035), .ZN(n2923) );
  inv0d1 U23 ( .I(n2969), .ZN(n3035) );
  nd04d0 U24 ( .A1(n1811), .A2(n1810), .A3(n1809), .A4(n1808), .ZN(n1812) );
  nd04d0 U25 ( .A1(n1799), .A2(n1798), .A3(n1797), .A4(n1796), .ZN(n1815) );
  nd04d0 U26 ( .A1(n1986), .A2(n1985), .A3(n1984), .A4(n1983), .ZN(n2001) );
  nd04d0 U27 ( .A1(n1992), .A2(n1991), .A3(n1990), .A4(n1989), .ZN(n2000) );
  nd04d0 U28 ( .A1(n1632), .A2(n1631), .A3(n1630), .A4(n1629), .ZN(n1648) );
  nd04d0 U29 ( .A1(n1980), .A2(n1979), .A3(n1978), .A4(n1977), .ZN(n2002) );
  nd04d0 U30 ( .A1(n1433), .A2(n1432), .A3(n1431), .A4(n1430), .ZN(n1434) );
  nd04d0 U31 ( .A1(n1462), .A2(n1461), .A3(n1460), .A4(n1459), .ZN(n1480) );
  nd04d0 U32 ( .A1(n1526), .A2(n1525), .A3(n1524), .A4(n1523), .ZN(n1542) );
  nd04d0 U33 ( .A1(n1476), .A2(n1475), .A3(n1474), .A4(n1473), .ZN(n1477) );
  nd04d0 U34 ( .A1(n1717), .A2(n1716), .A3(n1715), .A4(n1714), .ZN(n1734) );
  nd04d0 U35 ( .A1(n1320), .A2(n1319), .A3(n1318), .A4(n1317), .ZN(n1352) );
  nd04d0 U36 ( .A1(n1335), .A2(n1334), .A3(n1333), .A4(n1332), .ZN(n1350) );
  nd04d0 U37 ( .A1(n1920), .A2(n1919), .A3(n1918), .A4(n1917), .ZN(n1921) );
  nd04d0 U38 ( .A1(n1803), .A2(n1802), .A3(n1801), .A4(n1800), .ZN(n1814) );
  nd04d0 U39 ( .A1(n1730), .A2(n1729), .A3(n1728), .A4(n1727), .ZN(n1731) );
  nd04d0 U40 ( .A1(n1411), .A2(n1410), .A3(n1409), .A4(n1408), .ZN(n1412) );
  nd04d0 U41 ( .A1(n1348), .A2(n1347), .A3(n1346), .A4(n1345), .ZN(n1349) );
  nd04d0 U42 ( .A1(n1767), .A2(n1766), .A3(n1765), .A4(n1764), .ZN(n1773) );
  nd04d0 U43 ( .A1(n1467), .A2(n1466), .A3(n1465), .A4(n1464), .ZN(n1479) );
  nd04d0 U44 ( .A1(n1709), .A2(n1708), .A3(n1707), .A4(n1706), .ZN(n1710) );
  nd04d0 U45 ( .A1(n1701), .A2(n1700), .A3(n1699), .A4(n1698), .ZN(n1712) );
  nd04d0 U46 ( .A1(n1429), .A2(n1428), .A3(n1427), .A4(n1426), .ZN(n1435) );
  nd04d0 U47 ( .A1(n1998), .A2(n1997), .A3(n1996), .A4(n1995), .ZN(n1999) );
  nd04d0 U48 ( .A1(n1687), .A2(n1686), .A3(n1685), .A4(n1684), .ZN(n1688) );
  nd04d0 U49 ( .A1(n1891), .A2(n1890), .A3(n1889), .A4(n1888), .ZN(n1898) );
  nd04d0 U50 ( .A1(n1853), .A2(n1852), .A3(n1851), .A4(n1850), .ZN(n1854) );
  nd04d0 U51 ( .A1(n1849), .A2(n1848), .A3(n1847), .A4(n1846), .ZN(n1855) );
  nd04d0 U52 ( .A1(n1807), .A2(n1806), .A3(n1805), .A4(n1804), .ZN(n1813) );
  nd04d0 U53 ( .A1(n1845), .A2(n1844), .A3(n1843), .A4(n1842), .ZN(n1856) );
  nd04d0 U54 ( .A1(n1449), .A2(n1448), .A3(n1447), .A4(n1446), .ZN(n1455) );
  nd04d0 U55 ( .A1(n1832), .A2(n1831), .A3(n1830), .A4(n1829), .ZN(n1833) );
  nd04d0 U56 ( .A1(n1763), .A2(n1762), .A3(n1761), .A4(n1760), .ZN(n1774) );
  nd04d0 U57 ( .A1(n1841), .A2(n1840), .A3(n1839), .A4(n1838), .ZN(n1857) );
  nd04d0 U58 ( .A1(n1364), .A2(n1363), .A3(n1362), .A4(n1361), .ZN(n1370) );
  nd04d0 U59 ( .A1(n1445), .A2(n1444), .A3(n1443), .A4(n1442), .ZN(n1456) );
  nd04d0 U60 ( .A1(n1726), .A2(n1725), .A3(n1724), .A4(n1723), .ZN(n1732) );
  nd04d0 U61 ( .A1(n1329), .A2(n1328), .A3(n1327), .A4(n1326), .ZN(n1351) );
  nd04d0 U62 ( .A1(n1820), .A2(n1819), .A3(n1818), .A4(n1817), .ZN(n1836) );
  nd04d0 U63 ( .A1(n1356), .A2(n1355), .A3(n1354), .A4(n1353), .ZN(n1372) );
  nd04d0 U64 ( .A1(n1425), .A2(n1424), .A3(n1423), .A4(n1422), .ZN(n1436) );
  nd04d0 U65 ( .A1(n1828), .A2(n1827), .A3(n1826), .A4(n1825), .ZN(n1834) );
  nd04d0 U66 ( .A1(n1441), .A2(n1440), .A3(n1439), .A4(n1438), .ZN(n1457) );
  nd04d0 U67 ( .A1(n1360), .A2(n1359), .A3(n1358), .A4(n1357), .ZN(n1371) );
  nd04d0 U68 ( .A1(n1824), .A2(n1823), .A3(n1822), .A4(n1821), .ZN(n1835) );
  nd04d0 U69 ( .A1(n1421), .A2(n1420), .A3(n1419), .A4(n1418), .ZN(n1437) );
  nd04d0 U70 ( .A1(n1887), .A2(n1886), .A3(n1885), .A4(n1884), .ZN(n1899) );
  nd04d0 U71 ( .A1(n1705), .A2(n1704), .A3(n1703), .A4(n1702), .ZN(n1711) );
  nd04d0 U72 ( .A1(n1534), .A2(n1533), .A3(n1532), .A4(n1531), .ZN(n1540) );
  nd04d0 U73 ( .A1(n1611), .A2(n1610), .A3(n1609), .A4(n1608), .ZN(n1627) );
  nd04d0 U74 ( .A1(n1743), .A2(n1742), .A3(n1741), .A4(n1740), .ZN(n1754) );
  nd04d0 U75 ( .A1(n1572), .A2(n1571), .A3(n1570), .A4(n1569), .ZN(n1583) );
  nd04d0 U76 ( .A1(n1941), .A2(n1940), .A3(n1939), .A4(n1938), .ZN(n1949) );
  nd04d0 U77 ( .A1(n1513), .A2(n1512), .A3(n1511), .A4(n1510), .ZN(n1519) );
  nd04d0 U78 ( .A1(n1771), .A2(n1770), .A3(n1769), .A4(n1768), .ZN(n1772) );
  nd04d0 U79 ( .A1(n1568), .A2(n1567), .A3(n1566), .A4(n1565), .ZN(n1584) );
  nd04d0 U80 ( .A1(n1870), .A2(n1869), .A3(n1868), .A4(n1867), .ZN(n1876) );
  nd04d0 U81 ( .A1(n2037), .A2(n2036), .A3(n2035), .A4(n2034), .ZN(n2038) );
  nd04d0 U82 ( .A1(n1661), .A2(n1660), .A3(n1659), .A4(n1658), .ZN(n1667) );
  nd04d0 U83 ( .A1(n1739), .A2(n1738), .A3(n1737), .A4(n1736), .ZN(n1755) );
  nd04d0 U84 ( .A1(n1386), .A2(n1385), .A3(n1384), .A4(n1383), .ZN(n1393) );
  nd04d0 U85 ( .A1(n1589), .A2(n1588), .A3(n1587), .A4(n1586), .ZN(n1605) );
  nd04d0 U86 ( .A1(n1779), .A2(n1778), .A3(n1777), .A4(n1776), .ZN(n1795) );
  nd04d0 U87 ( .A1(n1747), .A2(n1746), .A3(n1745), .A4(n1744), .ZN(n1753) );
  nd04d0 U88 ( .A1(n1548), .A2(n1547), .A3(n1546), .A4(n1545), .ZN(n1564) );
  nd04d0 U89 ( .A1(n1675), .A2(n1674), .A3(n1673), .A4(n1672), .ZN(n1691) );
  nd04d0 U90 ( .A1(n1640), .A2(n1639), .A3(n1638), .A4(n1637), .ZN(n1646) );
  nd04d0 U91 ( .A1(n1957), .A2(n1956), .A3(n1955), .A4(n1954), .ZN(n1973) );
  nd04d0 U92 ( .A1(n1576), .A2(n1575), .A3(n1574), .A4(n1573), .ZN(n1582) );
  nd04d0 U93 ( .A1(n1615), .A2(n1614), .A3(n1613), .A4(n1612), .ZN(n1626) );
  nd04d0 U94 ( .A1(n1657), .A2(n1656), .A3(n1655), .A4(n1654), .ZN(n1668) );
  nd04d0 U95 ( .A1(n1947), .A2(n1946), .A3(n1945), .A4(n1944), .ZN(n1948) );
  nd04d0 U96 ( .A1(n1636), .A2(n1635), .A3(n1634), .A4(n1633), .ZN(n1647) );
  nd04d0 U97 ( .A1(n1560), .A2(n1559), .A3(n1558), .A4(n1557), .ZN(n1561) );
  nd04d0 U98 ( .A1(n1874), .A2(n1873), .A3(n1872), .A4(n1871), .ZN(n1875) );
  nd04d0 U99 ( .A1(n1623), .A2(n1622), .A3(n1621), .A4(n1620), .ZN(n1624) );
  nd04d0 U100 ( .A1(n1382), .A2(n1381), .A3(n1380), .A4(n1379), .ZN(n1394) );
  nd04d0 U101 ( .A1(n1783), .A2(n1782), .A3(n1781), .A4(n1780), .ZN(n1794) );
  nd04d0 U102 ( .A1(n1961), .A2(n1960), .A3(n1959), .A4(n1958), .ZN(n1972) );
  nd04d0 U103 ( .A1(n1911), .A2(n1910), .A3(n1909), .A4(n1908), .ZN(n1923) );
  nd04d0 U104 ( .A1(n2029), .A2(n2028), .A3(n2027), .A4(n2026), .ZN(n2039) );
  nd04d0 U105 ( .A1(n1751), .A2(n1750), .A3(n1749), .A4(n1748), .ZN(n1752) );
  nd04d0 U106 ( .A1(n1403), .A2(n1402), .A3(n1401), .A4(n1400), .ZN(n1414) );
  nd04d0 U107 ( .A1(n1376), .A2(n1375), .A3(n1374), .A4(n1373), .ZN(n1395) );
  nd04d0 U108 ( .A1(n1787), .A2(n1786), .A3(n1785), .A4(n1784), .ZN(n1793) );
  nd04d0 U109 ( .A1(n1679), .A2(n1678), .A3(n1677), .A4(n1676), .ZN(n1690) );
  nd04d0 U110 ( .A1(n1399), .A2(n1398), .A3(n1397), .A4(n1396), .ZN(n1415) );
  nd04d0 U111 ( .A1(n1915), .A2(n1914), .A3(n1913), .A4(n1912), .ZN(n1922) );
  nd04d0 U112 ( .A1(n1538), .A2(n1537), .A3(n1536), .A4(n1535), .ZN(n1539) );
  nd04d0 U113 ( .A1(n1492), .A2(n1491), .A3(n1490), .A4(n1489), .ZN(n1498) );
  nd04d0 U114 ( .A1(n1965), .A2(n1964), .A3(n1963), .A4(n1962), .ZN(n1971) );
  nd04d0 U115 ( .A1(n1517), .A2(n1516), .A3(n1515), .A4(n1514), .ZN(n1518) );
  nd04d0 U116 ( .A1(n1505), .A2(n1504), .A3(n1503), .A4(n1502), .ZN(n1521) );
  nd04d0 U117 ( .A1(n1930), .A2(n1929), .A3(n1928), .A4(n1927), .ZN(n1951) );
  nd04d0 U118 ( .A1(n1969), .A2(n1968), .A3(n1967), .A4(n1966), .ZN(n1970) );
  nd04d0 U119 ( .A1(n2010), .A2(n2009), .A3(n2008), .A4(n2007), .ZN(n2041) );
  nd04d0 U120 ( .A1(n1791), .A2(n1790), .A3(n1789), .A4(n1788), .ZN(n1792) );
  nd04d0 U121 ( .A1(n1601), .A2(n1600), .A3(n1599), .A4(n1598), .ZN(n1602) );
  nd04d0 U122 ( .A1(n1866), .A2(n1865), .A3(n1864), .A4(n1863), .ZN(n1877) );
  nd04d0 U123 ( .A1(n1556), .A2(n1555), .A3(n1554), .A4(n1553), .ZN(n1562) );
  nd04d0 U124 ( .A1(n1484), .A2(n1483), .A3(n1482), .A4(n1481), .ZN(n1500) );
  nd04d0 U125 ( .A1(n1862), .A2(n1861), .A3(n1860), .A4(n1859), .ZN(n1878) );
  nd04d0 U126 ( .A1(n1552), .A2(n1551), .A3(n1550), .A4(n1549), .ZN(n1563) );
  nd04d0 U127 ( .A1(n1496), .A2(n1495), .A3(n1494), .A4(n1493), .ZN(n1497) );
  nd04d0 U128 ( .A1(n1653), .A2(n1652), .A3(n1651), .A4(n1650), .ZN(n1669) );
  nd04d0 U129 ( .A1(n1896), .A2(n1895), .A3(n1894), .A4(n1893), .ZN(n1897) );
  nd04d0 U130 ( .A1(n1407), .A2(n1406), .A3(n1405), .A4(n1404), .ZN(n1413) );
  nd04d0 U131 ( .A1(n1683), .A2(n1682), .A3(n1681), .A4(n1680), .ZN(n1689) );
  nd04d0 U132 ( .A1(n1597), .A2(n1596), .A3(n1595), .A4(n1594), .ZN(n1603) );
  nd04d0 U133 ( .A1(n2019), .A2(n2018), .A3(n2017), .A4(n2016), .ZN(n2040) );
  nd04d0 U134 ( .A1(n1936), .A2(n1935), .A3(n1934), .A4(n1933), .ZN(n1950) );
  nd04d0 U135 ( .A1(n1619), .A2(n1618), .A3(n1617), .A4(n1616), .ZN(n1625) );
  nd04d0 U136 ( .A1(n1488), .A2(n1487), .A3(n1486), .A4(n1485), .ZN(n1499) );
  nd04d0 U137 ( .A1(n1883), .A2(n1882), .A3(n1881), .A4(n1880), .ZN(n1900) );
  nd04d0 U138 ( .A1(n1227), .A2(n1226), .A3(n1225), .A4(n1224), .ZN(n1235) );
  nd04d0 U139 ( .A1(n1221), .A2(n1220), .A3(n1219), .A4(n1218), .ZN(n1236) );
  nd04d0 U140 ( .A1(n657), .A2(n656), .A3(n655), .A4(n654), .ZN(n674) );
  nd04d0 U141 ( .A1(n824), .A2(n823), .A3(n822), .A4(n821), .ZN(n840) );
  nd04d0 U142 ( .A1(n678), .A2(n677), .A3(n676), .A4(n675), .ZN(n694) );
  nd04d0 U143 ( .A1(n1233), .A2(n1232), .A3(n1231), .A4(n1230), .ZN(n1234) );
  nd04d0 U144 ( .A1(n662), .A2(n661), .A3(n660), .A4(n659), .ZN(n673) );
  nd04d0 U145 ( .A1(n1001), .A2(n1000), .A3(n999), .A4(n998), .ZN(n1007) );
  nd04d0 U146 ( .A1(n1111), .A2(n1110), .A3(n1109), .A4(n1108), .ZN(n1112) );
  nd04d0 U147 ( .A1(n723), .A2(n722), .A3(n721), .A4(n720), .ZN(n734) );
  nd04d0 U148 ( .A1(n686), .A2(n685), .A3(n684), .A4(n683), .ZN(n692) );
  nd04d0 U149 ( .A1(n636), .A2(n635), .A3(n634), .A4(n633), .ZN(n652) );
  nd04d0 U150 ( .A1(n731), .A2(n730), .A3(n729), .A4(n728), .ZN(n732) );
  nd04d0 U151 ( .A1(n1189), .A2(n1188), .A3(n1187), .A4(n1186), .ZN(n1207) );
  nd04d0 U152 ( .A1(n1023), .A2(n1022), .A3(n1021), .A4(n1020), .ZN(n1029) );
  nd04d0 U153 ( .A1(n1214), .A2(n1213), .A3(n1212), .A4(n1211), .ZN(n1237) );
  nd04d0 U154 ( .A1(n997), .A2(n996), .A3(n995), .A4(n994), .ZN(n1008) );
  nd04d0 U155 ( .A1(n993), .A2(n992), .A3(n991), .A4(n990), .ZN(n1009) );
  nd04d0 U156 ( .A1(n832), .A2(n831), .A3(n830), .A4(n829), .ZN(n838) );
  nd04d0 U157 ( .A1(n1035), .A2(n1034), .A3(n1033), .A4(n1032), .ZN(n1051) );
  nd04d0 U158 ( .A1(n1039), .A2(n1038), .A3(n1037), .A4(n1036), .ZN(n1050) );
  nd04d0 U159 ( .A1(n1043), .A2(n1042), .A3(n1041), .A4(n1040), .ZN(n1049) );
  nd04d0 U160 ( .A1(n828), .A2(n827), .A3(n826), .A4(n825), .ZN(n839) );
  nd04d0 U161 ( .A1(n1089), .A2(n1088), .A3(n1087), .A4(n1086), .ZN(n1090) );
  nd04d0 U162 ( .A1(n875), .A2(n874), .A3(n873), .A4(n872), .ZN(n881) );
  nd04d0 U163 ( .A1(n1180), .A2(n1179), .A3(n1178), .A4(n1177), .ZN(n1181) );
  nd04d0 U164 ( .A1(n1085), .A2(n1084), .A3(n1083), .A4(n1082), .ZN(n1091) );
  nd04d0 U165 ( .A1(n1175), .A2(n1174), .A3(n1173), .A4(n1172), .ZN(n1182) );
  nd04d0 U166 ( .A1(n1081), .A2(n1080), .A3(n1079), .A4(n1078), .ZN(n1092) );
  nd04d0 U167 ( .A1(n1077), .A2(n1076), .A3(n1075), .A4(n1074), .ZN(n1093) );
  nd04d0 U168 ( .A1(n1170), .A2(n1169), .A3(n1168), .A4(n1167), .ZN(n1183) );
  nd04d0 U169 ( .A1(n1165), .A2(n1164), .A3(n1163), .A4(n1162), .ZN(n1184) );
  nd04d0 U170 ( .A1(n1098), .A2(n1097), .A3(n1096), .A4(n1095), .ZN(n1115) );
  nd04d0 U171 ( .A1(n1103), .A2(n1102), .A3(n1101), .A4(n1100), .ZN(n1114) );
  nd04d0 U172 ( .A1(n784), .A2(n783), .A3(n782), .A4(n781), .ZN(n800) );
  nd04d0 U173 ( .A1(n888), .A2(n887), .A3(n886), .A4(n885), .ZN(n905) );
  nd04d0 U174 ( .A1(n893), .A2(n892), .A3(n891), .A4(n890), .ZN(n904) );
  nd04d0 U175 ( .A1(n788), .A2(n787), .A3(n786), .A4(n785), .ZN(n799) );
  nd04d0 U176 ( .A1(n871), .A2(n870), .A3(n869), .A4(n868), .ZN(n882) );
  nd04d0 U177 ( .A1(n909), .A2(n908), .A3(n907), .A4(n906), .ZN(n925) );
  nd04d0 U178 ( .A1(n913), .A2(n912), .A3(n911), .A4(n910), .ZN(n924) );
  nd04d0 U179 ( .A1(n917), .A2(n916), .A3(n915), .A4(n914), .ZN(n923) );
  nd04d0 U180 ( .A1(n921), .A2(n920), .A3(n919), .A4(n918), .ZN(n922) );
  nd04d0 U181 ( .A1(n866), .A2(n865), .A3(n864), .A4(n863), .ZN(n883) );
  nd04d0 U182 ( .A1(n1055), .A2(n1054), .A3(n1053), .A4(n1052), .ZN(n1071) );
  nd04d0 U183 ( .A1(n1107), .A2(n1106), .A3(n1105), .A4(n1104), .ZN(n1113) );
  nd04d0 U184 ( .A1(n1059), .A2(n1058), .A3(n1057), .A4(n1056), .ZN(n1070) );
  nd04d0 U185 ( .A1(n594), .A2(n593), .A3(n592), .A4(n591), .ZN(n609) );
  nd04d0 U186 ( .A1(n942), .A2(n941), .A3(n940), .A4(n939), .ZN(n943) );
  nd04d0 U187 ( .A1(n792), .A2(n791), .A3(n790), .A4(n789), .ZN(n798) );
  nd04d0 U188 ( .A1(n711), .A2(n710), .A3(n709), .A4(n708), .ZN(n712) );
  nd04d0 U189 ( .A1(n707), .A2(n706), .A3(n705), .A4(n704), .ZN(n713) );
  nd04d0 U190 ( .A1(n587), .A2(n586), .A3(n585), .A4(n584), .ZN(n610) );
  nd04d0 U191 ( .A1(n703), .A2(n702), .A3(n701), .A4(n700), .ZN(n714) );
  nd04d0 U192 ( .A1(n698), .A2(n697), .A3(n696), .A4(n695), .ZN(n715) );
  nd04d0 U193 ( .A1(n938), .A2(n937), .A3(n936), .A4(n935), .ZN(n944) );
  nd04d0 U194 ( .A1(n577), .A2(n576), .A3(n575), .A4(n574), .ZN(n611) );
  nd04d0 U195 ( .A1(n934), .A2(n933), .A3(n932), .A4(n931), .ZN(n945) );
  nd04d0 U196 ( .A1(n1249), .A2(n1248), .A3(n1247), .A4(n1246), .ZN(n1267) );
  nd04d0 U197 ( .A1(n930), .A2(n929), .A3(n928), .A4(n927), .ZN(n946) );
  nd04d0 U198 ( .A1(n1063), .A2(n1062), .A3(n1061), .A4(n1060), .ZN(n1069) );
  nd04d0 U199 ( .A1(n1257), .A2(n1256), .A3(n1255), .A4(n1254), .ZN(n1266) );
  nd04d0 U200 ( .A1(n1264), .A2(n1263), .A3(n1262), .A4(n1261), .ZN(n1265) );
  nd04d0 U201 ( .A1(n1199), .A2(n1198), .A3(n1197), .A4(n1196), .ZN(n1205) );
  nd04d0 U202 ( .A1(n804), .A2(n803), .A3(n802), .A4(n801), .ZN(n820) );
  nd04d0 U203 ( .A1(n616), .A2(n615), .A3(n614), .A4(n613), .ZN(n632) );
  nd04d0 U204 ( .A1(n1133), .A2(n1132), .A3(n1131), .A4(n1130), .ZN(n1134) );
  nd04d0 U205 ( .A1(n748), .A2(n747), .A3(n746), .A4(n745), .ZN(n754) );
  nd04d0 U206 ( .A1(n770), .A2(n769), .A3(n768), .A4(n767), .ZN(n776) );
  nd04d0 U207 ( .A1(n744), .A2(n743), .A3(n742), .A4(n741), .ZN(n755) );
  nd04d0 U208 ( .A1(n644), .A2(n643), .A3(n642), .A4(n641), .ZN(n650) );
  nd04d0 U209 ( .A1(n1279), .A2(n1278), .A3(n1277), .A4(n1276), .ZN(n1306) );
  nd04d0 U210 ( .A1(n620), .A2(n619), .A3(n618), .A4(n617), .ZN(n631) );
  nd04d0 U211 ( .A1(n1286), .A2(n1285), .A3(n1284), .A4(n1283), .ZN(n1305) );
  nd04d0 U212 ( .A1(n740), .A2(n739), .A3(n738), .A4(n737), .ZN(n756) );
  nd04d0 U213 ( .A1(n666), .A2(n665), .A3(n664), .A4(n663), .ZN(n672) );
  nd04d0 U214 ( .A1(n1019), .A2(n1018), .A3(n1017), .A4(n1016), .ZN(n1030) );
  nd04d0 U215 ( .A1(n1293), .A2(n1292), .A3(n1291), .A4(n1290), .ZN(n1304) );
  nd04d0 U216 ( .A1(n954), .A2(n953), .A3(n952), .A4(n951), .ZN(n965) );
  nd04d0 U217 ( .A1(n1120), .A2(n1119), .A3(n1118), .A4(n1117), .ZN(n1137) );
  nd04d0 U218 ( .A1(n1129), .A2(n1128), .A3(n1127), .A4(n1126), .ZN(n1135) );
  nd04d0 U219 ( .A1(n978), .A2(n977), .A3(n976), .A4(n975), .ZN(n984) );
  nd04d0 U220 ( .A1(n624), .A2(n623), .A3(n622), .A4(n621), .ZN(n630) );
  nd04d0 U221 ( .A1(n1142), .A2(n1141), .A3(n1140), .A4(n1139), .ZN(n1160) );
  nd04d0 U222 ( .A1(n950), .A2(n949), .A3(n948), .A4(n947), .ZN(n966) );
  nd04d0 U223 ( .A1(n970), .A2(n969), .A3(n968), .A4(n967), .ZN(n986) );
  nd04d0 U224 ( .A1(n1125), .A2(n1124), .A3(n1123), .A4(n1122), .ZN(n1136) );
  nd04d0 U225 ( .A1(n1147), .A2(n1146), .A3(n1145), .A4(n1144), .ZN(n1159) );
  nd04d0 U226 ( .A1(n808), .A2(n807), .A3(n806), .A4(n805), .ZN(n819) );
  nd04d0 U227 ( .A1(n974), .A2(n973), .A3(n972), .A4(n971), .ZN(n985) );
  nd04d0 U228 ( .A1(n812), .A2(n811), .A3(n810), .A4(n809), .ZN(n818) );
  nd04d0 U229 ( .A1(n1152), .A2(n1151), .A3(n1150), .A4(n1149), .ZN(n1158) );
  nd04d0 U230 ( .A1(n719), .A2(n718), .A3(n717), .A4(n716), .ZN(n735) );
  nd04d0 U231 ( .A1(n846), .A2(n845), .A3(n844), .A4(n843), .ZN(n862) );
  nd04d0 U232 ( .A1(n958), .A2(n957), .A3(n956), .A4(n955), .ZN(n964) );
  nd04d0 U233 ( .A1(n1005), .A2(n1004), .A3(n1003), .A4(n1002), .ZN(n1006) );
  nd04d0 U234 ( .A1(n762), .A2(n761), .A3(n760), .A4(n759), .ZN(n778) );
  nd04d0 U235 ( .A1(n850), .A2(n849), .A3(n848), .A4(n847), .ZN(n861) );
  nd04d0 U236 ( .A1(n1015), .A2(n1014), .A3(n1013), .A4(n1012), .ZN(n1031) );
  nd04d0 U237 ( .A1(n640), .A2(n639), .A3(n638), .A4(n637), .ZN(n651) );
  nd04d0 U238 ( .A1(n766), .A2(n765), .A3(n764), .A4(n763), .ZN(n777) );
  nd04d0 U239 ( .A1(n854), .A2(n853), .A3(n852), .A4(n851), .ZN(n860) );
  nd04d0 U240 ( .A1(n392), .A2(n391), .A3(n390), .A4(n389), .ZN(n5935) );
  nd04d0 U241 ( .A1(n7007), .A2(n2371), .A3(n2370), .A4(n2369), .ZN(n2375) );
  nd04d0 U242 ( .A1(n379), .A2(n378), .A3(n377), .A4(n376), .ZN(n5932) );
  nd04d0 U243 ( .A1(n404), .A2(n403), .A3(n402), .A4(n401), .ZN(n5934) );
  nd04d0 U244 ( .A1(n325), .A2(n324), .A3(n323), .A4(n322), .ZN(n5931) );
  nd04d0 U245 ( .A1(n6503), .A2(n6502), .A3(n6501), .A4(n6500), .ZN(n6509) );
  nd04d0 U246 ( .A1(n6545), .A2(n6544), .A3(n6543), .A4(n6542), .ZN(n6546) );
  nd04d0 U247 ( .A1(n6532), .A2(n6531), .A3(n6530), .A4(n6529), .ZN(n6533) );
  nd04d0 U248 ( .A1(n6491), .A2(n6490), .A3(n6489), .A4(n6488), .ZN(n6497) );
  nd04d0 U249 ( .A1(n6507), .A2(n6506), .A3(n6505), .A4(n6504), .ZN(n6508) );
  nd04d0 U250 ( .A1(n6519), .A2(n6518), .A3(n6517), .A4(n6516), .ZN(n6520) );
  nd04d0 U251 ( .A1(n6527), .A2(n6526), .A3(n6525), .A4(n6524), .ZN(n6534) );
  nd04d0 U252 ( .A1(n4061), .A2(n4026), .A3(n4022), .A4(n3830), .ZN(n4079) );
  nd04d0 U253 ( .A1(n3829), .A2(n3828), .A3(n3827), .A4(n3826), .ZN(n5319) );
  nd04d0 U254 ( .A1(n3716), .A2(n3715), .A3(n3714), .A4(n3713), .ZN(n3731) );
  nd04d0 U255 ( .A1(n6122), .A2(n6121), .A3(n5323), .A4(n5322), .ZN(n6253) );
  nd04d0 U256 ( .A1(n6429), .A2(n6428), .A3(n6427), .A4(n6426), .ZN(n6430) );
  nd04d0 U257 ( .A1(n6425), .A2(n6424), .A3(n6423), .A4(n6422), .ZN(n6431) );
  nd04d0 U258 ( .A1(n6442), .A2(n6441), .A3(n6440), .A4(n6439), .ZN(n6443) );
  nd04d0 U259 ( .A1(n6437), .A2(n6436), .A3(n6435), .A4(n6434), .ZN(n6444) );
  nd04d0 U260 ( .A1(n6454), .A2(n6453), .A3(n6452), .A4(n6451), .ZN(n6455) );
  nd04d0 U261 ( .A1(n6450), .A2(n6449), .A3(n6448), .A4(n6447), .ZN(n6456) );
  nd04d0 U262 ( .A1(n6464), .A2(n6463), .A3(n6462), .A4(n6461), .ZN(n6471) );
  nd04d0 U263 ( .A1(n6483), .A2(n6482), .A3(n6481), .A4(n6480), .ZN(n6484) );
  nd04d0 U264 ( .A1(n6479), .A2(n6478), .A3(n6477), .A4(n6476), .ZN(n6485) );
  nd04d0 U265 ( .A1(n6495), .A2(n6494), .A3(n6493), .A4(n6492), .ZN(n6496) );
  nd04d0 U266 ( .A1(n6632), .A2(n6631), .A3(n6630), .A4(n6629), .ZN(n6633) );
  nd04d0 U267 ( .A1(n6627), .A2(n6626), .A3(n6625), .A4(n6624), .ZN(n6634) );
  nd04d0 U268 ( .A1(n6645), .A2(n6644), .A3(n6643), .A4(n6642), .ZN(n6646) );
  nd04d0 U269 ( .A1(n6641), .A2(n6640), .A3(n6639), .A4(n6638), .ZN(n6647) );
  nd04d0 U270 ( .A1(n6656), .A2(n6655), .A3(n6654), .A4(n6653), .ZN(n6662) );
  nd04d0 U271 ( .A1(n6676), .A2(n6675), .A3(n6674), .A4(n6673), .ZN(n6677) );
  nd04d0 U272 ( .A1(n6670), .A2(n6669), .A3(n6668), .A4(n6667), .ZN(n6678) );
  nd04d0 U273 ( .A1(n6689), .A2(n6688), .A3(n6687), .A4(n6686), .ZN(n6690) );
  nd04d0 U274 ( .A1(n6685), .A2(n6684), .A3(n6683), .A4(n6682), .ZN(n6691) );
  nd04d0 U275 ( .A1(n6704), .A2(n6703), .A3(n6702), .A4(n6701), .ZN(n6705) );
  nd04d0 U276 ( .A1(n6700), .A2(n6699), .A3(n6698), .A4(n6697), .ZN(n6706) );
  nd04d0 U277 ( .A1(n6717), .A2(n6716), .A3(n6715), .A4(n6714), .ZN(n6718) );
  nd04d0 U278 ( .A1(n6713), .A2(n6712), .A3(n6711), .A4(n6710), .ZN(n6719) );
  nd04d0 U279 ( .A1(n6733), .A2(n6732), .A3(n6731), .A4(n6730), .ZN(n6734) );
  nd04d0 U280 ( .A1(n6727), .A2(n6726), .A3(n6725), .A4(n6724), .ZN(n6735) );
  nd04d0 U281 ( .A1(n6748), .A2(n6747), .A3(n6746), .A4(n6745), .ZN(n6749) );
  nd04d0 U282 ( .A1(n6744), .A2(n6743), .A3(n6742), .A4(n6741), .ZN(n6750) );
  nd04d0 U283 ( .A1(n6762), .A2(n6761), .A3(n6760), .A4(n6759), .ZN(n6763) );
  nd04d0 U284 ( .A1(n6758), .A2(n6757), .A3(n6756), .A4(n6755), .ZN(n6764) );
  nd04d0 U285 ( .A1(n6776), .A2(n6775), .A3(n6774), .A4(n6773), .ZN(n6777) );
  nd04d0 U286 ( .A1(n6795), .A2(n6794), .A3(n6793), .A4(n6792), .ZN(n6796) );
  nd04d0 U287 ( .A1(n6788), .A2(n6787), .A3(n6786), .A4(n6785), .ZN(n6797) );
  nd04d0 U288 ( .A1(n7106), .A2(n7105), .A3(n7104), .A4(n7103), .ZN(n7108) );
  nd04d0 U289 ( .A1(n7101), .A2(n7100), .A3(n7099), .A4(n7098), .ZN(n7109) );
  nd04d0 U290 ( .A1(n6607), .A2(n6606), .A3(n6605), .A4(n6604), .ZN(n6608) );
  nd04d0 U291 ( .A1(n6570), .A2(n6569), .A3(n6568), .A4(n6567), .ZN(n6571) );
  nd04d0 U292 ( .A1(n6603), .A2(n6602), .A3(n6601), .A4(n6600), .ZN(n6609) );
  nd04d0 U293 ( .A1(n6578), .A2(n6577), .A3(n6576), .A4(n6575), .ZN(n6584) );
  nd04d0 U294 ( .A1(n6619), .A2(n6618), .A3(n6617), .A4(n6616), .ZN(n6620) );
  nd04d0 U295 ( .A1(n6594), .A2(n6593), .A3(n6592), .A4(n6591), .ZN(n6595) );
  nd04d0 U296 ( .A1(n6558), .A2(n6557), .A3(n6556), .A4(n6555), .ZN(n6559) );
  nd04d0 U297 ( .A1(n6553), .A2(n6552), .A3(n6551), .A4(n6550), .ZN(n6560) );
  nd04d0 U298 ( .A1(n6615), .A2(n6614), .A3(n6613), .A4(n6612), .ZN(n6621) );
  nd04d0 U299 ( .A1(n6590), .A2(n6589), .A3(n6588), .A4(n6587), .ZN(n6596) );
  nd04d0 U300 ( .A1(n6541), .A2(n6540), .A3(n6539), .A4(n6538), .ZN(n6547) );
  nd04d0 U301 ( .A1(n6515), .A2(n6514), .A3(n6513), .A4(n6512), .ZN(n6521) );
  nd04d0 U302 ( .A1(n6582), .A2(n6581), .A3(n6580), .A4(n6579), .ZN(n6583) );
  nd04d0 U303 ( .A1(n3044), .A2(n3000), .A3(n353), .A4(n2631), .ZN(n218) );
  nd04d0 U304 ( .A1(n3815), .A2(n3814), .A3(n3813), .A4(n3812), .ZN(n3816) );
  nd04d0 U305 ( .A1(n281), .A2(n264), .A3(n263), .A4(n262), .ZN(n271) );
  nd04d0 U306 ( .A1(n2364), .A2(
        \IBusCachedPlugin_cache/_zz_when_InstructionCache_l342 ), .A3(n2363), 
        .A4(n2425), .ZN(n2365) );
  nd04d0 U307 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n3795), .ZN(n3809) );
  nd04d0 U308 ( .A1(HazardSimplePlugin_writeBackBuffer_valid), .A2(n238), .A3(
        n237), .A4(n236), .ZN(n239) );
  nd04d0 U309 ( .A1(HazardSimplePlugin_writeBackBuffer_valid), .A2(n260), .A3(
        n259), .A4(n258), .ZN(n277) );
  nd04d0 U310 ( .A1(n288), .A2(n287), .A3(n2247), .A4(n286), .ZN(n289) );
  nd04d0 U311 ( .A1(n2623), .A2(n2618), .A3(n174), .A4(n2622), .ZN(n183) );
  nr02d0 U312 ( .A1(n1312), .A2(n1314), .ZN(n1322) );
  nr02d0 U313 ( .A1(n1312), .A2(n1307), .ZN(n1315) );
  nd02d0 U314 ( .A1(n1316), .A2(n1315), .ZN(n1342) );
  nd02d0 U315 ( .A1(n1321), .A2(n1323), .ZN(n1343) );
  nd02d0 U316 ( .A1(n1322), .A2(n1323), .ZN(n1330) );
  nd02d0 U317 ( .A1(n1316), .A2(n1324), .ZN(n1337) );
  nd02d0 U318 ( .A1(n1316), .A2(n1322), .ZN(n1339) );
  nd02d0 U319 ( .A1(n1311), .A2(n1310), .ZN(n1344) );
  nd02d0 U320 ( .A1(n1309), .A2(n1310), .ZN(n1341) );
  nd02d0 U321 ( .A1(n1315), .A2(n1323), .ZN(n1336) );
  nd02d0 U322 ( .A1(n1308), .A2(n1309), .ZN(n1340) );
  nd02d0 U323 ( .A1(n1324), .A2(n1323), .ZN(n1338) );
  nd02d0 U324 ( .A1(n1311), .A2(n1308), .ZN(n1331) );
  nd02d0 U325 ( .A1(n1316), .A2(n1321), .ZN(n1325) );
  nd02d0 U326 ( .A1(n573), .A2(n582), .ZN(n595) );
  nd02d0 U327 ( .A1(n580), .A2(n573), .ZN(n598) );
  nd02d0 U328 ( .A1(n580), .A2(n583), .ZN(n589) );
  nd02d0 U329 ( .A1(n580), .A2(n570), .ZN(n601) );
  nd02d0 U330 ( .A1(n572), .A2(n568), .ZN(n597) );
  nd02d0 U331 ( .A1(n581), .A2(n582), .ZN(n588) );
  nd02d0 U332 ( .A1(n571), .A2(n569), .ZN(n590) );
  nd02d0 U333 ( .A1(n583), .A2(n582), .ZN(n602) );
  nd02d0 U334 ( .A1(n569), .A2(n568), .ZN(n603) );
  nd02d0 U335 ( .A1(n580), .A2(n581), .ZN(n596) );
  nd02d0 U336 ( .A1(n572), .A2(n571), .ZN(n600) );
  nd02d0 U337 ( .A1(n570), .A2(n582), .ZN(n599) );
  ad01d0 U338 ( .A(n3016), .B(n3002), .CI(n3001), .CO(n354), .S(n3004) );
  ad01d0 U339 ( .A(n563), .B(n355), .CI(n354), .CO(n2976), .S(n356) );
  ad01d0 U340 ( .A(n2990), .B(n2977), .CI(n2976), .CO(n2962), .S(n2978) );
  ad01d0 U341 ( .A(n2965), .B(n2963), .CI(n2962), .CO(n2948), .S(n2964) );
  ad01d0 U342 ( .A(n2951), .B(n2949), .CI(n2948), .CO(n2928), .S(n2950) );
  ad01d0 U343 ( .A(n2931), .B(n2929), .CI(n2928), .CO(n2911), .S(n2930) );
  ad01d0 U344 ( .A(n2914), .B(n2912), .CI(n2911), .CO(n2895), .S(n2913) );
  ad01d0 U345 ( .A(n2899), .B(n2896), .CI(n2895), .CO(n2882), .S(n2898) );
  ad01d0 U346 ( .A(n2885), .B(n2883), .CI(n2882), .CO(n2864), .S(n2884) );
  ad01d0 U347 ( .A(n2873), .B(n2865), .CI(n2864), .CO(n339), .S(n2866) );
  ad01d0 U348 ( .A(n2869), .B(n340), .CI(n339), .CO(n369), .S(n312) );
  ad01d0 U349 ( .A(n2291), .B(n370), .CI(n369), .CO(n2849), .S(n371) );
  ad01d0 U350 ( .A(n2863), .B(n2850), .CI(n2849), .CO(n394), .S(n2851) );
  ad01d0 U351 ( .A(n2848), .B(n395), .CI(n394), .CO(n382), .S(n396) );
  ad01d0 U352 ( .A(n2282), .B(n383), .CI(n382), .CO(n2830), .S(n384) );
  ad01d0 U353 ( .A(n2838), .B(n2831), .CI(n2830), .CO(n2815), .S(n2832) );
  ad01d0 U354 ( .A(n2835), .B(n2816), .CI(n2815), .CO(n2801), .S(n2817) );
  ad01d0 U355 ( .A(n2812), .B(n2802), .CI(n2801), .CO(n2787), .S(n2803) );
  ad01d0 U356 ( .A(n2805), .B(n2788), .CI(n2787), .CO(n2771), .S(n2789) );
  ad01d0 U357 ( .A(n2782), .B(n2772), .CI(n2771), .CO(n2118), .S(n2773) );
  ad01d0 U358 ( .A(n2775), .B(n2119), .CI(n2118), .CO(n2756), .S(n341) );
  ad01d0 U359 ( .A(n2760), .B(n2757), .CI(n2756), .CO(n2736), .S(n2758) );
  ad01d0 U360 ( .A(n2728), .B(n2726), .CI(n2725), .CO(n2708), .S(n2727) );
  ad01d0 U361 ( .A(n2711), .B(n2699), .CI(n2698), .CO(n2679), .S(n2700) );
  ad01d0 U362 ( .A(n2694), .B(n2680), .CI(n2679), .CO(n2667), .S(n2681) );
  ad01d0 U363 ( .A(n2670), .B(n2668), .CI(n2667), .CO(n2650), .S(n2669) );
  ad01d0 U364 ( .A(n2659), .B(n2651), .CI(n2650), .CO(n2120), .S(n2652) );
  ad01d0 U365 ( .A(n3039), .B(n311), .CI(n310), .CO(n3001), .S(n219) );
  ad01d0 U366 ( .A(n2644), .B(n220), .CI(execute_SRC_USE_SUB_LESS), .CO(n310), 
        .S(n221) );
  nd03d0 U367 ( .A1(n3316), .A2(n3315), .A3(n3314), .ZN(n3498) );
  nd03d0 U368 ( .A1(n2614), .A2(n2613), .A3(n2612), .ZN(n2098) );
  ad01d0 U369 ( .A(n2740), .B(n2737), .CI(n2736), .CO(n2725), .S(n2738) );
  ad01d0 U370 ( .A(n2713), .B(n2709), .CI(n2708), .CO(n2698), .S(n2710) );
  nd03d0 U371 ( .A1(n3683), .A2(n3695), .A3(n3690), .ZN(n2354) );
  nd02d0 U372 ( .A1(n212), .A2(n211), .ZN(n2988) );
  nd02d0 U373 ( .A1(n2601), .A2(n2597), .ZN(n336) );
  nd02d0 U374 ( .A1(execute_arbitration_isValid), .A2(execute_IS_CSR), .ZN(
        n562) );
  nd02d0 U375 ( .A1(n222), .A2(n2289), .ZN(n6998) );
  ad01d0 U376 ( .A(n6414), .B(n6413), .CI(n6412), .CO(n6408), .S(n6415) );
  ad01d0 U377 ( .A(n6410), .B(n6409), .CI(n6408), .CO(n6404), .S(n6411) );
  ad01d0 U378 ( .A(n6406), .B(n6405), .CI(n6404), .CO(n6400), .S(n6407) );
  ad01d0 U379 ( .A(n6402), .B(n6401), .CI(n6400), .CO(n6397), .S(n6403) );
  ad01d0 U380 ( .A(_zz__zz_execute_SRC2_3[5]), .B(n6398), .CI(n6397), .CO(
        n6394), .S(n6399) );
  ad01d0 U381 ( .A(_zz__zz_execute_SRC2_3[6]), .B(n6395), .CI(n6394), .CO(
        n6391), .S(n6396) );
  ad01d0 U382 ( .A(_zz__zz_execute_SRC2_3[7]), .B(n6392), .CI(n6391), .CO(
        n6388), .S(n6393) );
  ad01d0 U383 ( .A(_zz__zz_execute_SRC2_3[8]), .B(n6389), .CI(n6388), .CO(
        n6385), .S(n6390) );
  ad01d0 U384 ( .A(_zz__zz_execute_SRC2_3[9]), .B(n6386), .CI(n6385), .CO(
        n6382), .S(n6387) );
  ad01d0 U385 ( .A(_zz__zz_execute_SRC2_3[10]), .B(n6383), .CI(n6382), .CO(
        n6378), .S(n6384) );
  ad01d0 U386 ( .A(n6380), .B(n6379), .CI(n6378), .CO(n6374), .S(n6381) );
  ad01d0 U387 ( .A(n6376), .B(n6375), .CI(n6374), .CO(n6370), .S(n6377) );
  ad01d0 U388 ( .A(n6372), .B(n6371), .CI(n6370), .CO(n6366), .S(n6373) );
  ad01d0 U389 ( .A(n6368), .B(n6367), .CI(n6366), .CO(n6362), .S(n6369) );
  ad01d0 U390 ( .A(n6364), .B(n6363), .CI(n6362), .CO(n6358), .S(n6365) );
  ad01d0 U391 ( .A(n6360), .B(n6359), .CI(n6358), .CO(n6354), .S(n6361) );
  ad01d0 U392 ( .A(n6356), .B(n6355), .CI(n6354), .CO(n6350), .S(n6357) );
  ad01d0 U393 ( .A(n6352), .B(n6351), .CI(n6350), .CO(n6346), .S(n6353) );
  ad01d0 U394 ( .A(n6348), .B(n6347), .CI(n6346), .CO(n6342), .S(n6349) );
  ad01d0 U395 ( .A(n6344), .B(n6343), .CI(n6342), .CO(n6339), .S(n6345) );
  ad01d0 U396 ( .A(n6340), .B(n6343), .CI(n6339), .CO(n6336), .S(n6341) );
  ad01d0 U397 ( .A(n6337), .B(_zz__zz_execute_SRC2_3[11]), .CI(n6336), .CO(
        n6333), .S(n6338) );
  ad01d0 U398 ( .A(n6334), .B(_zz__zz_execute_SRC2_3[11]), .CI(n6333), .CO(
        n6330), .S(n6335) );
  ad01d0 U399 ( .A(n6331), .B(_zz__zz_execute_SRC2_3[11]), .CI(n6330), .CO(
        n6327), .S(n6332) );
  ad01d0 U400 ( .A(n6328), .B(_zz__zz_execute_SRC2_3[11]), .CI(n6327), .CO(
        n6324), .S(n6329) );
  ad01d0 U401 ( .A(n6325), .B(_zz__zz_execute_SRC2_3[11]), .CI(n6324), .CO(
        n6321), .S(n6326) );
  ad01d0 U402 ( .A(n6322), .B(n6343), .CI(n6321), .CO(n6318), .S(n6323) );
  ad01d0 U403 ( .A(n6319), .B(n6343), .CI(n6318), .CO(n6315), .S(n6320) );
  ad01d0 U404 ( .A(n6316), .B(n6343), .CI(n6315), .CO(n6312), .S(n6317) );
  ad01d0 U405 ( .A(n6313), .B(n6343), .CI(n6312), .CO(n6309), .S(n6314) );
  nd02d0 U406 ( .A1(execute_arbitration_isValid), .A2(execute_DO_EBREAK), .ZN(
        n2474) );
  nd02d0 U407 ( .A1(execute_CsrPlugin_csr_833), .A2(n3566), .ZN(n3666) );
  nd03d0 U408 ( .A1(n2555), .A2(n3045), .A3(n2591), .ZN(n2571) );
  nr03d0 U409 ( .A1(n562), .A2(n3238), .A3(n2551), .ZN(n3566) );
  nd03d0 U410 ( .A1(n2547), .A2(n2616), .A3(n2610), .ZN(n2546) );
  nd03d0 U411 ( .A1(n2403), .A2(n6740), .A3(n7121), .ZN(n2240) );
  nd03d0 U412 ( .A1(n2358), .A2(n2360), .A3(n2357), .ZN(n2242) );
  nd03d0 U413 ( .A1(n2358), .A2(n3049), .A3(n2357), .ZN(n2373) );
  nd03d0 U414 ( .A1(n3040), .A2(n2282), .A3(n388), .ZN(n389) );
  nd03d0 U415 ( .A1(n2310), .A2(n2309), .A3(n2308), .ZN(n2926) );
  nd02d0 U416 ( .A1(n2749), .A2(n562), .ZN(n3033) );
  nd03d0 U417 ( .A1(n431), .A2(n430), .A3(n429), .ZN(n6112) );
  nd03d0 U418 ( .A1(n451), .A2(n450), .A3(n449), .ZN(n6106) );
  nd03d0 U419 ( .A1(n547), .A2(n546), .A3(n545), .ZN(n6105) );
  nd03d0 U420 ( .A1(n497), .A2(n496), .A3(n495), .ZN(n6104) );
  nd03d0 U421 ( .A1(n462), .A2(n461), .A3(n460), .ZN(n6097) );
  nd03d0 U422 ( .A1(n482), .A2(n481), .A3(n480), .ZN(n6095) );
  nd03d0 U423 ( .A1(n467), .A2(n466), .A3(n465), .ZN(n6094) );
  nd03d0 U424 ( .A1(n2232), .A2(n7121), .A3(n2231), .ZN(n2230) );
  nd03d0 U425 ( .A1(n2744), .A2(n2743), .A3(n2742), .ZN(n2745) );
  nd03d0 U426 ( .A1(n2716), .A2(n2715), .A3(n2714), .ZN(n2717) );
  nd03d0 U427 ( .A1(n519), .A2(n518), .A3(n517), .ZN(n6089) );
  nd03d0 U428 ( .A1(n364), .A2(n363), .A3(n362), .ZN(n5922) );
  inv0d0 U429 ( .I(decode_INSTRUCTION[18]), .ZN(n173) );
  inv0d0 U430 ( .I(decode_INSTRUCTION[15]), .ZN(n174) );
  nd02d2 U431 ( .A1(execute_SRC1_CTRL[0]), .A2(n2601), .ZN(n302) );
  inv0d1 U432 ( .I(n6666), .ZN(n2266) );
  nd02d4 U433 ( .A1(n7007), .A2(n7006), .ZN(n7077) );
  nr02d4 U434 ( .A1(n7006), .A2(n3719), .ZN(n6651) );
  nr02d4 U435 ( .A1(n7006), .A2(n3712), .ZN(n6672) );
  inv0d1 U436 ( .I(n3056), .ZN(n3058) );
  inv0d2 U437 ( .I(iBus_rsp_payload_data[25]), .ZN(n3178) );
  inv0d2 U438 ( .I(n6301), .ZN(n6290) );
  nr03d1 U439 ( .A1(n2403), .A2(n2394), .A3(n2405), .ZN(n416) );
  inv0d1 U440 ( .I(n6996), .ZN(n7116) );
  inv0d1 U441 ( .I(decode_INSTRUCTION_24), .ZN(n2613) );
  inv0d2 U442 ( .I(n3287), .ZN(n3499) );
  inv0d2 U443 ( .I(n2476), .ZN(n2526) );
  inv0d2 U444 ( .I(execute_CsrPlugin_csr_833), .ZN(n2541) );
  inv0d2 U445 ( .I(iBus_rsp_payload_data[31]), .ZN(n3166) );
  inv0d2 U446 ( .I(n6908), .ZN(n6893) );
  inv0d2 U447 ( .I(n2856), .ZN(n2996) );
  inv0d4 U448 ( .I(n2594), .ZN(n2117) );
  inv0d1 U449 ( .I(decode_INSTRUCTION_22), .ZN(n2615) );
  inv0d1 U450 ( .I(decode_INSTRUCTION[19]), .ZN(n2618) );
  inv0d1 U451 ( .I(execute_ALU_BITWISE_CTRL[1]), .ZN(n6681) );
  nd02d2 U452 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3263), .ZN(n3342)
         );
  nd02d2 U453 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3265), .ZN(n3344)
         );
  nr02d0 U454 ( .A1(n3709), .A2(n3708), .ZN(n3711) );
  nr02d0 U455 ( .A1(n3705), .A2(n3709), .ZN(n3722) );
  nd04d0 U456 ( .A1(n269), .A2(n268), .A3(n267), .A4(n266), .ZN(n270) );
  nd04d0 U457 ( .A1(n3769), .A2(n3768), .A3(n3767), .A4(n3766), .ZN(n3770) );
  nr02d0 U458 ( .A1(n1313), .A2(n1307), .ZN(n1321) );
  nr02d0 U459 ( .A1(n3016), .A2(n3015), .ZN(n3007) );
  nr02d0 U460 ( .A1(n7006), .A2(n3718), .ZN(n6528) );
  nr02d0 U461 ( .A1(n7005), .A2(n3718), .ZN(n6460) );
  nr04d0 U462 ( .A1(n3773), .A2(n3772), .A3(n3771), .A4(n3770), .ZN(n3774) );
  nr02d0 U463 ( .A1(n2483), .A2(n2484), .ZN(n2479) );
  nr02d0 U464 ( .A1(n1331), .A2(n1338), .ZN(n1463) );
  nr02d0 U465 ( .A1(n590), .A2(n601), .ZN(n612) );
  nd04d0 U466 ( .A1(n3433), .A2(n232), .A3(n231), .A4(n230), .ZN(n240) );
  nr02d0 U467 ( .A1(n2671), .A2(n2653), .ZN(n2654) );
  nr02d0 U468 ( .A1(n6306), .A2(n6305), .ZN(n6308) );
  nd04d0 U469 ( .A1(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[0] ), .A2(
        n3807), .A3(n3806), .A4(n3805), .ZN(n3808) );
  nd03d0 U470 ( .A1(n3776), .A2(n3775), .A3(n3774), .ZN(n3778) );
  nr02d0 U471 ( .A1(n1344), .A2(n1342), .ZN(n2005) );
  nr02d0 U472 ( .A1(n1341), .A2(n1338), .ZN(n1697) );
  nr02d0 U473 ( .A1(n597), .A2(n596), .ZN(n699) );
  nr02d0 U474 ( .A1(n600), .A2(n598), .ZN(n1185) );
  nr02d0 U475 ( .A1(n589), .A2(n603), .ZN(n780) );
  nr02d0 U476 ( .A1(n603), .A2(n588), .ZN(n1216) );
  nr02d0 U477 ( .A1(n1340), .A2(n1339), .ZN(n1472) );
  nr02d0 U478 ( .A1(n590), .A2(n595), .ZN(n736) );
  nr02d0 U479 ( .A1(n590), .A2(n588), .ZN(n1161) );
  nr02d0 U480 ( .A1(n1340), .A2(n1338), .ZN(n1378) );
  nr02d0 U481 ( .A1(n603), .A2(n598), .ZN(n989) );
  nr02d0 U482 ( .A1(n597), .A2(n599), .ZN(n987) );
  nr02d0 U483 ( .A1(n601), .A2(n603), .ZN(n758) );
  nd03d0 U484 ( .A1(n3309), .A2(n3315), .A3(n3314), .ZN(n3489) );
  nd02d0 U485 ( .A1(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[2] ), 
        .A2(n3159), .ZN(n3147) );
  nd12d0 U486 ( .A1(n2051), .A2(n2050), .ZN(n2053) );
  nd03d0 U487 ( .A1(n2761), .A2(n2760), .A3(n2759), .ZN(n2762) );
  nr02d0 U488 ( .A1(n2728), .A2(n2722), .ZN(n3749) );
  nr03d0 U489 ( .A1(n2682), .A2(n2666), .A3(n2961), .ZN(n2673) );
  nr03d0 U490 ( .A1(n2975), .A2(n2981), .A3(n2961), .ZN(n2968) );
  nr02d0 U491 ( .A1(n2198), .A2(n2214), .ZN(n2216) );
  nd04d0 U492 ( .A1(n6771), .A2(n6770), .A3(n6769), .A4(n6768), .ZN(n6778) );
  nd04d0 U493 ( .A1(n6660), .A2(n6659), .A3(n6658), .A4(n6657), .ZN(n6661) );
  nd04d0 U494 ( .A1(n6566), .A2(n6565), .A3(n6564), .A4(n6563), .ZN(n6572) );
  nd04d0 U495 ( .A1(n6469), .A2(n6468), .A3(n6467), .A4(n6466), .ZN(n6470) );
  nd04d0 U496 ( .A1(n6251), .A2(n6250), .A3(n6249), .A4(n6248), .ZN(n6252) );
  nd04d0 U497 ( .A1(n3729), .A2(n3728), .A3(n3727), .A4(n3726), .ZN(n3730) );
  nr02d0 U498 ( .A1(n2554), .A2(n2575), .ZN(n2361) );
  nr02d0 U499 ( .A1(n2111), .A2(n6291), .ZN(n2951) );
  nd03d0 U500 ( .A1(n2298), .A2(n2297), .A3(n2296), .ZN(n2871) );
  nr03d0 U501 ( .A1(n2268), .A2(n2775), .A3(n6919), .ZN(n2269) );
  nr02d0 U502 ( .A1(n2051), .A2(n558), .ZN(n2190) );
  nr03d0 U503 ( .A1(n2198), .A2(n2137), .A3(n2136), .ZN(n2150) );
  nd03d0 U504 ( .A1(n3433), .A2(n3432), .A3(n3431), .ZN(n3497) );
  nr02d0 U505 ( .A1(n3444), .A2(n3392), .ZN(n3370) );
  nr02d0 U506 ( .A1(n3317), .A2(n3449), .ZN(n3296) );
  nr02d0 U507 ( .A1(n2054), .A2(n2053), .ZN(n2368) );
  nr02d0 U508 ( .A1(n3158), .A2(n3147), .ZN(n3148) );
  nr02d0 U509 ( .A1(n3121), .A2(n3147), .ZN(n3102) );
  nr02d0 U510 ( .A1(n3049), .A2(n2214), .ZN(n2399) );
  nd04d0 U511 ( .A1(n352), .A2(n351), .A3(n350), .A4(n349), .ZN(n564) );
  nd12d0 U512 ( .A1(n304), .A2(n303), .ZN(n308) );
  nr02d0 U513 ( .A1(n295), .A2(n2242), .ZN(n561) );
  nd04d0 U514 ( .A1(n727), .A2(n726), .A3(n725), .A4(n724), .ZN(n733) );
  nd04d0 U515 ( .A1(n1644), .A2(n1643), .A3(n1642), .A4(n1641), .ZN(n1645) );
  nd04d0 U516 ( .A1(n1509), .A2(n1508), .A3(n1507), .A4(n1506), .ZN(n1520) );
  nd04d0 U517 ( .A1(n836), .A2(n835), .A3(n834), .A4(n833), .ZN(n837) );
  nd04d0 U518 ( .A1(n1696), .A2(n1695), .A3(n1694), .A4(n1693), .ZN(n1713) );
  nr03d0 U519 ( .A1(n3672), .A2(n2345), .A3(reset), .ZN(n2351) );
  nd02d1 U520 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3277), .ZN(n3465)
         );
  nd04d0 U521 ( .A1(n1156), .A2(n1155), .A3(n1154), .A4(n1153), .ZN(n1157) );
  nd04d0 U522 ( .A1(n1368), .A2(n1367), .A3(n1366), .A4(n1365), .ZN(n1369) );
  nd04d0 U523 ( .A1(n982), .A2(n981), .A3(n980), .A4(n979), .ZN(n983) );
  nd04d0 U524 ( .A1(n1722), .A2(n1721), .A3(n1720), .A4(n1719), .ZN(n1733) );
  nd04d0 U525 ( .A1(n1047), .A2(n1046), .A3(n1045), .A4(n1044), .ZN(n1048) );
  nr02d0 U526 ( .A1(CsrPlugin_mstatus_MPP[0]), .A2(n2342), .ZN(n2341) );
  nd04d0 U527 ( .A1(n1907), .A2(n1906), .A3(n1905), .A4(n1904), .ZN(n1924) );
  nd04d0 U528 ( .A1(n858), .A2(n857), .A3(n856), .A4(n855), .ZN(n859) );
  nd04d0 U529 ( .A1(n1203), .A2(n1202), .A3(n1201), .A4(n1200), .ZN(n1204) );
  nd04d0 U530 ( .A1(n1194), .A2(n1193), .A3(n1192), .A4(n1191), .ZN(n1206) );
  nd04d0 U531 ( .A1(n1243), .A2(n1242), .A3(n1241), .A4(n1240), .ZN(n1268) );
  nd04d0 U532 ( .A1(n1027), .A2(n1026), .A3(n1025), .A4(n1024), .ZN(n1028) );
  nd02d1 U533 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3268), .ZN(n3458)
         );
  nd04d0 U534 ( .A1(n796), .A2(n795), .A3(n794), .A4(n793), .ZN(n797) );
  nd04d0 U535 ( .A1(n1665), .A2(n1664), .A3(n1663), .A4(n1662), .ZN(n1666) );
  nd04d0 U536 ( .A1(n1302), .A2(n1301), .A3(n1300), .A4(n1299), .ZN(n1303) );
  nd04d0 U537 ( .A1(n1471), .A2(n1470), .A3(n1469), .A4(n1468), .ZN(n1478) );
  nd04d0 U538 ( .A1(n962), .A2(n961), .A3(n960), .A4(n959), .ZN(n963) );
  nd04d0 U539 ( .A1(n1593), .A2(n1592), .A3(n1591), .A4(n1590), .ZN(n1604) );
  nd04d0 U540 ( .A1(n879), .A2(n878), .A3(n877), .A4(n876), .ZN(n880) );
  nd04d0 U541 ( .A1(n1530), .A2(n1529), .A3(n1528), .A4(n1527), .ZN(n1541) );
  nd04d0 U542 ( .A1(n1067), .A2(n1066), .A3(n1065), .A4(n1064), .ZN(n1068) );
  nd04d0 U543 ( .A1(n1759), .A2(n1758), .A3(n1757), .A4(n1756), .ZN(n1775) );
  nd04d0 U544 ( .A1(n816), .A2(n815), .A3(n814), .A4(n813), .ZN(n817) );
  nd04d0 U545 ( .A1(n901), .A2(n900), .A3(n899), .A4(n898), .ZN(n902) );
  nd04d0 U546 ( .A1(n897), .A2(n896), .A3(n895), .A4(n894), .ZN(n903) );
  nd04d0 U547 ( .A1(n690), .A2(n689), .A3(n688), .A4(n687), .ZN(n691) );
  nd04d0 U548 ( .A1(n682), .A2(n681), .A3(n680), .A4(n679), .ZN(n693) );
  nd04d0 U549 ( .A1(n648), .A2(n647), .A3(n646), .A4(n645), .ZN(n649) );
  nd04d0 U550 ( .A1(n670), .A2(n669), .A3(n668), .A4(n667), .ZN(n671) );
  nd04d0 U551 ( .A1(n628), .A2(n627), .A3(n626), .A4(n625), .ZN(n629) );
  nd04d0 U552 ( .A1(n1453), .A2(n1452), .A3(n1451), .A4(n1450), .ZN(n1454) );
  nd04d0 U553 ( .A1(n752), .A2(n751), .A3(n750), .A4(n749), .ZN(n753) );
  nd04d0 U554 ( .A1(n1580), .A2(n1579), .A3(n1578), .A4(n1577), .ZN(n1581) );
  nd04d0 U555 ( .A1(n607), .A2(n606), .A3(n605), .A4(n604), .ZN(n608) );
  nd04d0 U556 ( .A1(n1391), .A2(n1390), .A3(n1389), .A4(n1388), .ZN(n1392) );
  nd04d0 U557 ( .A1(n774), .A2(n773), .A3(n772), .A4(n771), .ZN(n775) );
  nd02d1 U558 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3285), .ZN(n3473)
         );
  nd04d0 U559 ( .A1(n2589), .A2(n2616), .A3(n2617), .A4(n2610), .ZN(n2550) );
  nr03d0 U560 ( .A1(n3238), .A2(n2610), .A3(n2549), .ZN(n2540) );
  nd03d0 U561 ( .A1(n2403), .A2(n6996), .A3(n7121), .ZN(n2239) );
  nr02d0 U562 ( .A1(CsrPlugin_exceptionPendings_0), .A2(n285), .ZN(n2054) );
  nr04d0 U563 ( .A1(n2732), .A2(n2731), .A3(n2730), .A4(n2729), .ZN(n2735) );
  nr02d0 U564 ( .A1(n299), .A2(n2640), .ZN(n3697) );
  nr02d0 U565 ( .A1(n6740), .A2(n6781), .ZN(n3981) );
  nr02d0 U566 ( .A1(n3060), .A2(n293), .ZN(n6086) );
  nd03d0 U567 ( .A1(n457), .A2(n456), .A3(n455), .ZN(n6113) );
  nd03d0 U568 ( .A1(n524), .A2(n523), .A3(n522), .ZN(n6111) );
  nd03d0 U569 ( .A1(n502), .A2(n501), .A3(n500), .ZN(n6110) );
  nd03d0 U570 ( .A1(n426), .A2(n425), .A3(n424), .ZN(n6109) );
  nd03d0 U571 ( .A1(n446), .A2(n445), .A3(n444), .ZN(n6108) );
  nd03d0 U572 ( .A1(n530), .A2(n529), .A3(n528), .ZN(n6103) );
  nd03d0 U573 ( .A1(n487), .A2(n486), .A3(n485), .ZN(n6102) );
  nd03d0 U574 ( .A1(n472), .A2(n471), .A3(n470), .ZN(n6101) );
  nd03d0 U575 ( .A1(n514), .A2(n513), .A3(n512), .ZN(n6100) );
  nd03d0 U576 ( .A1(n477), .A2(n476), .A3(n475), .ZN(n6099) );
  nd03d0 U577 ( .A1(n492), .A2(n491), .A3(n490), .ZN(n6098) );
  nd03d0 U578 ( .A1(n410), .A2(n409), .A3(n408), .ZN(n6096) );
  nd03d0 U579 ( .A1(n415), .A2(n414), .A3(n413), .ZN(n6093) );
  nd03d0 U580 ( .A1(n436), .A2(n435), .A3(n434), .ZN(n6092) );
  nd03d0 U581 ( .A1(n537), .A2(n536), .A3(n535), .ZN(n6091) );
  nd03d0 U582 ( .A1(n421), .A2(n420), .A3(n419), .ZN(n6090) );
  nr02d0 U583 ( .A1(n2412), .A2(n248), .ZN(N1771) );
  nd03d0 U584 ( .A1(n210), .A2(n558), .A3(n2193), .ZN(n6208) );
  nr03d0 U585 ( .A1(n2412), .A2(DebugPlugin_godmode), .A3(n3250), .ZN(N1792)
         );
  nr02d0 U586 ( .A1(n2412), .A2(n2219), .ZN(N1840) );
  nd04d0 U587 ( .A1(n2427), .A2(n175), .A3(n179), .A4(n2226), .ZN(N2076) );
  nd03d0 U588 ( .A1(n441), .A2(n440), .A3(n439), .ZN(n6107) );
  nd03d0 U589 ( .A1(n348), .A2(n347), .A3(n346), .ZN(n5941) );
  nd03d0 U590 ( .A1(n509), .A2(n508), .A3(n507), .ZN(n6088) );
  nd03d0 U591 ( .A1(n292), .A2(n291), .A3(n290), .ZN(N2210) );
  inv0d1 U592 ( .I(reset), .ZN(n7121) );
  nr02d0 U593 ( .A1(memory_arbitration_isValid), .A2(lastStageIsValid), .ZN(
        n2427) );
  nr02d0 U594 ( .A1(IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid), 
        .A2(_zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1), .ZN(n175)
         );
  inv0d0 U595 ( .I(execute_arbitration_isValid), .ZN(n179) );
  inv0d0 U596 ( .I(switch_Fetcher_l362[2]), .ZN(n2234) );
  nd02d0 U597 ( .A1(switch_Fetcher_l362[1]), .A2(n2234), .ZN(n2226) );
  inv0d0 U598 ( .I(n7121), .ZN(n2412) );
  inv0d1 U599 ( .I(CsrPlugin_exceptionPendings_3), .ZN(n3250) );
  nd02d0 U600 ( .A1(lastStageIsValid), .A2(writeBack_REGFILE_WRITE_VALID), 
        .ZN(n248) );
  inv0d0 U601 ( .I(dBusWishbone_WE), .ZN(n6782) );
  aoi31d1 U602 ( .B1(n7265), .B2(dBusWishbone_ACK), .B3(n6782), .A(
        memory_MEMORY_STORE), .ZN(n176) );
  nd03d0 U603 ( .A1(memory_MEMORY_ENABLE), .A2(memory_arbitration_isValid), 
        .A3(n176), .ZN(n7117) );
  buffd1 U604 ( .I(n7117), .Z(n6926) );
  buffd1 U605 ( .I(n6926), .Z(n7113) );
  inv0d1 U606 ( .I(n7113), .ZN(n6889) );
  nd02d0 U607 ( .A1(memory_arbitration_isValid), .A2(memory_BRANCH_DO), .ZN(
        n2137) );
  inv0d0 U608 ( .I(memory_BRANCH_CALC[1]), .ZN(n2136) );
  nd03d0 U609 ( .A1(memory_MEMORY_ENABLE), .A2(memory_arbitration_isValid), 
        .A3(memory_ALIGNEMENT_FAULT), .ZN(n2135) );
  oai21d1 U610 ( .B1(n2137), .B2(n2136), .A(n2135), .ZN(n2241) );
  nr02d0 U611 ( .A1(n2241), .A2(CsrPlugin_exceptionPendings_2), .ZN(n2362) );
  inv0d0 U612 ( .I(lastStageIsValid), .ZN(n2046) );
  nr13d1 U613 ( .A1(writeBack_ENV_CTRL[0]), .A2(writeBack_ENV_CTRL[1]), .A3(
        n2046), .ZN(n405) );
  inv0d0 U614 ( .I(CsrPlugin_hadException), .ZN(n3673) );
  inv0d0 U615 ( .I(DebugPlugin_haltIt), .ZN(n2435) );
  inv0d0 U616 ( .I(DebugPlugin_stepIt), .ZN(n2422) );
  nd03d0 U617 ( .A1(CsrPlugin_interrupt_valid), .A2(n2435), .A3(n2422), .ZN(
        n295) );
  inv0d0 U618 ( .I(n295), .ZN(n273) );
  inv0d0 U619 ( .I(n3673), .ZN(n3671) );
  inv0d1 U620 ( .I(CsrPlugin_exceptionPendings_3), .ZN(n3245) );
  nr04d0 U621 ( .A1(n3671), .A2(CsrPlugin_exceptionPendings_3), .A3(
        CsrPlugin_exceptionPendings_2), .A4(CsrPlugin_exceptionPendings_1), 
        .ZN(n177) );
  nd03d0 U622 ( .A1(n273), .A2(CsrPlugin_pipelineLiberator_pcValids_2), .A3(
        n177), .ZN(n2534) );
  nd02d0 U623 ( .A1(n3673), .A2(n2534), .ZN(n3672) );
  nr02d0 U624 ( .A1(n405), .A2(n3672), .ZN(n2403) );
  inv0d0 U625 ( .I(n2403), .ZN(n2367) );
  nr04d0 U626 ( .A1(n6889), .A2(reset), .A3(n2362), .A4(n2367), .ZN(N1784) );
  buffd1 U627 ( .I(n7265), .Z(dBusWishbone_CYC) );
  inv0d0 U628 ( .I(\IBusCachedPlugin_cache/lineLoader_valid ), .ZN(n2413) );
  nr03d0 U629 ( .A1(iBusWishbone_ADR[0]), .A2(iBusWishbone_ADR[1]), .A3(
        iBusWishbone_ADR[2]), .ZN(n178) );
  oai21d1 U630 ( .B1(\IBusCachedPlugin_cache/lineLoader_cmdSent ), .B2(n2413), 
        .A(n178), .ZN(when_InstructionCache_l239) );
  inv0d0 U631 ( .I(iBusWishbone_ADR[3]), .ZN(\iBusWishbone_ADR[3]_BAR ) );
  inv0d0 U632 ( .I(execute_ENV_CTRL[1]), .ZN(n6802) );
  nr03d0 U633 ( .A1(execute_ENV_CTRL[0]), .A2(n6802), .A3(n179), .ZN(n2051) );
  inv0d0 U634 ( .I(n2241), .ZN(n209) );
  nd02d0 U635 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[6]), .A2(
        _zz_decode_LEGAL_INSTRUCTION_1[5]), .ZN(n207) );
  inv0d0 U636 ( .I(_zz_decode_LEGAL_INSTRUCTION_1[4]), .ZN(n2553) );
  nd02d0 U637 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[2]), .A2(n2553), .ZN(n206)
         );
  inv0d0 U638 ( .I(_zz_decode_LEGAL_INSTRUCTION_1[2]), .ZN(n3047) );
  nr02d0 U639 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[6]), .A2(n3047), .ZN(n2595)
         );
  nr03d0 U640 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[4]), .A2(
        _zz_decode_LEGAL_INSTRUCTION_1_13), .A3(
        \_zz_decode_LEGAL_INSTRUCTION_7[14] ), .ZN(n186) );
  inv0d0 U641 ( .I(_zz_decode_LEGAL_INSTRUCTION_1[5]), .ZN(n2630) );
  inv0d0 U642 ( .I(_zz_decode_LEGAL_INSTRUCTION_1[3]), .ZN(n2575) );
  aoi31d1 U643 ( .B1(n2595), .B2(n186), .B3(n2630), .A(n2575), .ZN(n205) );
  inv0d0 U644 ( .I(_zz_decode_LEGAL_INSTRUCTION_7_12), .ZN(n2554) );
  inv0d0 U645 ( .I(_zz_decode_LEGAL_INSTRUCTION_1_13), .ZN(n2072) );
  nd02d0 U646 ( .A1(n2554), .A2(n2072), .ZN(n2578) );
  inv0d0 U647 ( .I(n2578), .ZN(n2434) );
  nr02d0 U648 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[4]), .A2(
        \_zz_decode_LEGAL_INSTRUCTION_7[14] ), .ZN(n203) );
  inv0d0 U649 ( .I(n207), .ZN(n202) );
  inv0d0 U650 ( .I(decode_INSTRUCTION_10), .ZN(n2628) );
  inv0d0 U651 ( .I(decode_INSTRUCTION_11), .ZN(n2627) );
  nd02d0 U652 ( .A1(n2628), .A2(n2627), .ZN(n180) );
  nr04d0 U653 ( .A1(decode_INSTRUCTION_7), .A2(decode_INSTRUCTION_8), .A3(
        decode_INSTRUCTION_9), .A4(n180), .ZN(n2580) );
  inv0d0 U654 ( .I(_zz_decode_LEGAL_INSTRUCTION_13[26]), .ZN(n2610) );
  inv0d0 U655 ( .I(\_zz_decode_LEGAL_INSTRUCTION_7[14] ), .ZN(n2625) );
  nd04d0 U656 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[4]), .A2(n2580), .A3(n2610), 
        .A4(n2625), .ZN(n189) );
  inv0d0 U657 ( .I(_zz_decode_LEGAL_INSTRUCTION_13[28]), .ZN(n2606) );
  nr02d0 U658 ( .A1(decode_INSTRUCTION_22), .A2(n2606), .ZN(n2559) );
  aoi31d1 U659 ( .B1(\_zz__zz_decode_ENV_CTRL_2_1[20] ), .B2(
        _zz_decode_LEGAL_INSTRUCTION_1[6]), .B3(
        _zz_decode_LEGAL_INSTRUCTION_13[28]), .A(n2615), .ZN(n181) );
  nr04d0 U660 ( .A1(decode_INSTRUCTION_21), .A2(
        _zz_decode_LEGAL_INSTRUCTION_13[29]), .A3(n2559), .A4(n181), .ZN(n185)
         );
  inv0d1 U661 ( .I(decode_INSTRUCTION_21), .ZN(n2616) );
  nd02d0 U662 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[6]), .A2(
        _zz_decode_LEGAL_INSTRUCTION_13[28]), .ZN(n182) );
  nr04d0 U663 ( .A1(\_zz__zz_decode_ENV_CTRL_2_1[20] ), .A2(
        decode_INSTRUCTION_22), .A3(n2616), .A4(n182), .ZN(n184) );
  inv0d0 U664 ( .I(decode_INSTRUCTION_23), .ZN(n2614) );
  inv0d0 U665 ( .I(_zz_decode_LEGAL_INSTRUCTION_13[25]), .ZN(n2612) );
  nr04d0 U666 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13[27]), .A2(
        decode_INSTRUCTION_30), .A3(_zz_decode_LEGAL_INSTRUCTION_13_31), .A4(
        n2098), .ZN(n2543) );
  inv0d0 U667 ( .I(decode_INSTRUCTION[16]), .ZN(n2623) );
  inv0d0 U668 ( .I(decode_INSTRUCTION[15]), .ZN(n2624) );
  inv0d0 U669 ( .I(decode_INSTRUCTION[17]), .ZN(n2622) );
  nr02d0 U670 ( .A1(decode_INSTRUCTION[18]), .A2(n183), .ZN(n2552) );
  oai211d1 U671 ( .C1(n185), .C2(n184), .A(n2543), .B(n2552), .ZN(n188) );
  inv0d0 U672 ( .I(n186), .ZN(n187) );
  nd03d0 U673 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[4]), .A2(
        _zz_decode_LEGAL_INSTRUCTION_1[6]), .A3(n2578), .ZN(n2563) );
  oai211d1 U674 ( .C1(n189), .C2(n188), .A(n187), .B(n2563), .ZN(n190) );
  aoi31d1 U675 ( .B1(_zz_decode_LEGAL_INSTRUCTION_1[6]), .B2(
        \_zz_decode_LEGAL_INSTRUCTION_7[14] ), .B3(n2553), .A(n190), .ZN(n200)
         );
  nd02d0 U676 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[5]), .A2(n3047), .ZN(n2556)
         );
  nr02d0 U677 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13[27]), .A2(
        _zz_decode_LEGAL_INSTRUCTION_13_31), .ZN(n198) );
  nr02d0 U678 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[2]), .A2(
        \_zz_decode_LEGAL_INSTRUCTION_7[14] ), .ZN(n2585) );
  inv0d0 U679 ( .I(decode_INSTRUCTION_30), .ZN(n2605) );
  aoi31d1 U680 ( .B1(_zz_decode_LEGAL_INSTRUCTION_7_12), .B2(
        \_zz_decode_LEGAL_INSTRUCTION_7[14] ), .B3(n2072), .A(n2605), .ZN(n191) );
  aoi211d1 U681 ( .C1(_zz_decode_LEGAL_INSTRUCTION_1[5]), .C2(
        _zz_decode_LEGAL_INSTRUCTION_13[25]), .A(n191), .B(n2553), .ZN(n192)
         );
  aoi31d1 U682 ( .B1(n2585), .B2(n2434), .B3(n2612), .A(n192), .ZN(n193) );
  nr04d0 U683 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13[26]), .A2(
        _zz_decode_LEGAL_INSTRUCTION_13[28]), .A3(
        _zz_decode_LEGAL_INSTRUCTION_13[29]), .A4(n193), .ZN(n197) );
  inv0d0 U684 ( .I(n206), .ZN(n2598) );
  oai211d1 U685 ( .C1(_zz_decode_LEGAL_INSTRUCTION_1[4]), .C2(
        _zz_decode_LEGAL_INSTRUCTION_1_13), .A(
        _zz_decode_LEGAL_INSTRUCTION_7_12), .B(n3047), .ZN(n194) );
  aoi22d1 U686 ( .A1(n203), .A2(n2554), .B1(n2556), .B2(n194), .ZN(n195) );
  nd02d0 U687 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[4]), .A2(
        _zz_decode_LEGAL_INSTRUCTION_1_13), .ZN(n2586) );
  oai22d1 U688 ( .A1(n2598), .A2(n195), .B1(_zz_decode_LEGAL_INSTRUCTION_1[5]), 
        .B2(n2586), .ZN(n196) );
  inv0d0 U689 ( .I(_zz_decode_LEGAL_INSTRUCTION_1[6]), .ZN(n2577) );
  aon211d1 U690 ( .C1(n198), .C2(n197), .B(n196), .A(n2577), .ZN(n199) );
  oai211d1 U691 ( .C1(n200), .C2(n2556), .A(n2575), .B(n199), .ZN(n201) );
  aoi31d1 U692 ( .B1(n2434), .B2(n203), .B3(n202), .A(n201), .ZN(n204) );
  oan211d1 U693 ( .C1(n207), .C2(n206), .B(n205), .A(n204), .ZN(n208) );
  inv0d0 U694 ( .I(\IBusCachedPlugin_cache/decodeStage_hit_valid ), .ZN(n3817)
         );
  inv0d0 U695 ( .I(IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid), 
        .ZN(n2359) );
  oai21d1 U696 ( .B1(n3817), .B2(n2359), .A(n2226), .ZN(n2360) );
  inv0d0 U697 ( .I(n2360), .ZN(n2426) );
  aoi31d1 U698 ( .B1(_zz_decode_LEGAL_INSTRUCTION_1[0]), .B2(
        _zz_decode_LEGAL_INSTRUCTION_1[1]), .B3(n208), .A(n2426), .ZN(n285) );
  inv0d0 U699 ( .I(n285), .ZN(n2357) );
  nd02d0 U700 ( .A1(n209), .A2(n2357), .ZN(n2134) );
  nr02d0 U701 ( .A1(n2051), .A2(n2134), .ZN(n2181) );
  buffd1 U702 ( .I(n2181), .Z(n2204) );
  aoi22d1 U703 ( .A1(memory_MEMORY_STORE), .A2(n2198), .B1(n2204), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_code[1]), .ZN(n210) );
  nd02d0 U704 ( .A1(n285), .A2(n209), .ZN(n558) );
  nd02d0 U705 ( .A1(n2051), .A2(n209), .ZN(n2189) );
  buffd1 U706 ( .I(n2189), .Z(n2193) );
  inv0d0 U707 ( .I(execute_SHIFT_CTRL[1]), .ZN(n2572) );
  inv0d0 U708 ( .I(execute_SHIFT_CTRL[0]), .ZN(n2570) );
  inv0d0 U709 ( .I(execute_SRC2_CTRL[0]), .ZN(n2581) );
  nr02d0 U710 ( .A1(execute_SRC2_CTRL[1]), .A2(n2581), .ZN(n304) );
  inv0d0 U711 ( .I(execute_SRC2_CTRL[1]), .ZN(n2584) );
  nr02d1 U712 ( .A1(n2581), .A2(n2584), .ZN(n2105) );
  buffd1 U713 ( .I(n2105), .Z(n2113) );
  aoi22d1 U714 ( .A1(n304), .A2(_zz__zz_execute_BranchPlugin_branch_src2_3), 
        .B1(n2113), .B2(execute_PC[4]), .ZN(n212) );
  nr02d0 U715 ( .A1(execute_SRC2_CTRL[0]), .A2(execute_SRC2_CTRL[1]), .ZN(
        n2103) );
  buffd1 U716 ( .I(n2103), .Z(n2114) );
  nr02d0 U717 ( .A1(execute_SRC2_CTRL[0]), .A2(n2584), .ZN(n217) );
  aoi22d1 U718 ( .A1(n2114), .A2(execute_RS2[4]), .B1(n217), .B2(
        _zz__zz_execute_SRC2_3[4]), .ZN(n211) );
  aoi222d1 U719 ( .A1(n2114), .A2(execute_RS2[1]), .B1(
        _zz__zz_execute_SRC2_3[1]), .B2(n217), .C1(n304), .C2(
        _zz__zz_execute_BranchPlugin_branch_src2_0), .ZN(n3044) );
  inv0d0 U720 ( .I(n217), .ZN(n303) );
  inv0d0 U721 ( .I(_zz__zz_execute_SRC2_3[2]), .ZN(n6722) );
  buffd1 U722 ( .I(n2103), .Z(n2109) );
  aoi22d1 U723 ( .A1(n2109), .A2(execute_RS2[2]), .B1(n2113), .B2(
        execute_PC[2]), .ZN(n213) );
  oai21d1 U724 ( .B1(n303), .B2(n6722), .A(n213), .ZN(n214) );
  aoi21d1 U725 ( .B1(n304), .B2(_zz__zz_execute_BranchPlugin_branch_src2_1), 
        .A(n214), .ZN(n3000) );
  inv0d0 U726 ( .I(_zz__zz_execute_SRC2_3[3]), .ZN(n6709) );
  aoi22d1 U727 ( .A1(n2109), .A2(execute_RS2[3]), .B1(n304), .B2(
        _zz__zz_execute_BranchPlugin_branch_src2_2), .ZN(n215) );
  oai21d1 U728 ( .B1(n303), .B2(n6709), .A(n215), .ZN(n216) );
  aoi21d1 U729 ( .B1(n2113), .B2(execute_PC[3]), .A(n216), .ZN(n353) );
  aoi222d1 U730 ( .A1(n2114), .A2(execute_RS2[0]), .B1(n217), .B2(
        _zz__zz_execute_SRC2_3[0]), .C1(n304), .C2(
        _zz__zz_execute_BranchPlugin_branch_src2[10]), .ZN(n2631) );
  oai21d1 U731 ( .B1(n2988), .B2(n218), .A(execute_arbitration_isValid), .ZN(
        n315) );
  aoi21d1 U732 ( .B1(n2572), .B2(n2570), .A(n315), .ZN(n300) );
  inv0d0 U733 ( .I(execute_LightShifterPlugin_isActive), .ZN(n3679) );
  inv0d0 U734 ( .I(n3044), .ZN(n3038) );
  oai22d1 U735 ( .A1(n3679), .A2(execute_LightShifterPlugin_amplitudeReg[1]), 
        .B1(n3038), .B2(execute_LightShifterPlugin_isActive), .ZN(n3680) );
  inv0d0 U736 ( .I(n3680), .ZN(n3686) );
  inv0d0 U737 ( .I(execute_LightShifterPlugin_amplitudeReg[2]), .ZN(n3688) );
  aoi22d1 U738 ( .A1(execute_LightShifterPlugin_isActive), .A2(n3688), .B1(
        n3000), .B2(n3679), .ZN(n3685) );
  nr02d0 U739 ( .A1(n3686), .A2(n3685), .ZN(n3683) );
  aoi22d1 U740 ( .A1(execute_LightShifterPlugin_isActive), .A2(
        execute_LightShifterPlugin_amplitudeReg[4]), .B1(n2988), .B2(n3679), 
        .ZN(n3695) );
  inv0d0 U741 ( .I(n353), .ZN(n361) );
  aoi22d1 U742 ( .A1(execute_LightShifterPlugin_isActive), .A2(
        execute_LightShifterPlugin_amplitudeReg[3]), .B1(n361), .B2(n3679), 
        .ZN(n3690) );
  buffd1 U743 ( .I(n7117), .Z(n6997) );
  buffd1 U744 ( .I(n6997), .Z(n6996) );
  nd02d1 U745 ( .A1(n6996), .A2(n2474), .ZN(n299) );
  buffd1 U746 ( .I(n7265), .Z(n6977) );
  inv0d0 U747 ( .I(n6977), .ZN(n6993) );
  inv0d0 U748 ( .I(execute_SRC1_CTRL[1]), .ZN(n2601) );
  inv0d0 U749 ( .I(execute_SRC1_CTRL[0]), .ZN(n2597) );
  buffd3 U750 ( .I(n336), .Z(n2111) );
  inv0d0 U751 ( .I(execute_RS1[1]), .ZN(n6304) );
  nd02d0 U752 ( .A1(execute_SRC1_CTRL[1]), .A2(execute_SRC1_CTRL[0]), .ZN(n309) );
  inv0d0 U753 ( .I(_zz__zz_execute_SRC1_1[1]), .ZN(n6275) );
  oai22d1 U754 ( .A1(n2111), .A2(n6304), .B1(n309), .B2(n6275), .ZN(n3039) );
  inv0d1 U755 ( .I(execute_SRC_USE_SUB_LESS), .ZN(n2110) );
  inv0d1 U756 ( .I(execute_SRC_USE_SUB_LESS), .ZN(n2594) );
  aoi22d1 U757 ( .A1(n3044), .A2(n2110), .B1(n2117), .B2(n3038), .ZN(n311) );
  inv0d0 U758 ( .I(execute_RS1[0]), .ZN(n6306) );
  inv0d0 U759 ( .I(_zz__zz_execute_SRC1_1[0]), .ZN(n6277) );
  oai22d1 U760 ( .A1(n2111), .A2(n6306), .B1(n309), .B2(n6277), .ZN(n2644) );
  inv0d0 U761 ( .I(n2631), .ZN(n3678) );
  aoi22d1 U762 ( .A1(n2631), .A2(n2594), .B1(n2117), .B2(n3678), .ZN(n220) );
  inv0d1 U763 ( .I(execute_SRC2_FORCE_ZERO), .ZN(n3003) );
  aoi22d1 U764 ( .A1(execute_SRC2_FORCE_ZERO), .A2(n3039), .B1(n219), .B2(
        n3003), .ZN(n6981) );
  inv0d0 U765 ( .I(_zz__zz_execute_BranchPlugin_branch_src2[12]), .ZN(n6919)
         );
  inv0d1 U766 ( .I(execute_SRC2_FORCE_ZERO), .ZN(n2897) );
  aoi22d1 U767 ( .A1(execute_SRC2_FORCE_ZERO), .A2(n2644), .B1(n221), .B2(
        n2897), .ZN(n6994) );
  inv0d0 U768 ( .I(_zz__zz_execute_BranchPlugin_branch_src2[12]), .ZN(n6666)
         );
  nr02d0 U769 ( .A1(n2266), .A2(execute_ALU_BITWISE_CTRL[1]), .ZN(n556) );
  oan211d1 U770 ( .C1(n6981), .C2(n6919), .B(n6994), .A(n556), .ZN(n222) );
  nd02d1 U771 ( .A1(_zz__zz_execute_BranchPlugin_branch_src2[12]), .A2(
        execute_ALU_BITWISE_CTRL[1]), .ZN(n2331) );
  buffd1 U772 ( .I(n2331), .Z(n2289) );
  nd03d0 U773 ( .A1(execute_arbitration_isValid), .A2(execute_MEMORY_ENABLE), 
        .A3(n6998), .ZN(n2213) );
  oai22d1 U774 ( .A1(n2427), .A2(n562), .B1(n6993), .B2(n2213), .ZN(n223) );
  aor211d1 U775 ( .C1(n300), .C2(n2354), .A(n299), .B(n223), .Z(n3235) );
  buffd1 U776 ( .I(n3235), .Z(n3243) );
  buffd1 U777 ( .I(n3243), .Z(n2621) );
  inv0d1 U778 ( .I(n2621), .ZN(n2589) );
  inv0d0 U779 ( .I(memory_ENV_CTRL[1]), .ZN(n6803) );
  aoi31d1 U780 ( .B1(memory_arbitration_isValid), .B2(memory_ENV_CTRL[0]), 
        .B3(n6803), .A(n405), .ZN(n284) );
  nr02d0 U781 ( .A1(switch_Fetcher_l362[0]), .A2(n2226), .ZN(n2225) );
  aoi31d1 U782 ( .B1(execute_arbitration_isValid), .B2(execute_ENV_CTRL[0]), 
        .B3(n6802), .A(n2225), .ZN(n283) );
  aoi21d1 U783 ( .B1(_zz_decode_LEGAL_INSTRUCTION_1[6]), .B2(
        _zz_decode_LEGAL_INSTRUCTION_1[4]), .A(n2556), .ZN(n281) );
  oai221d1 U784 ( .B1(n2615), .B2(memory_INSTRUCTION[9]), .C1(n2614), .C2(
        memory_INSTRUCTION[10]), .A(n224), .ZN(n242) );
  inv0d0 U785 ( .I(\_zz__zz_decode_ENV_CTRL_2_1[20] ), .ZN(n2617) );
  oai22d1 U786 ( .A1(n2617), .A2(memory_INSTRUCTION[7]), .B1(n2616), .B2(
        memory_INSTRUCTION[8]), .ZN(n225) );
  aoi221d1 U787 ( .B1(n2617), .B2(memory_INSTRUCTION[7]), .C1(
        memory_INSTRUCTION[8]), .C2(n2616), .A(n225), .ZN(n227) );
  inv0d0 U788 ( .I(memory_INSTRUCTION[11]), .ZN(n6695) );
  aoi22d1 U789 ( .A1(decode_INSTRUCTION_24), .A2(n6695), .B1(
        memory_INSTRUCTION[11]), .B2(n2613), .ZN(n226) );
  nd04d0 U790 ( .A1(memory_REGFILE_WRITE_VALID), .A2(
        memory_arbitration_isValid), .A3(n227), .A4(n226), .ZN(n241) );
  inv0d0 U791 ( .I(n248), .ZN(n3433) );
  oai22d1 U792 ( .A1(_zz_lastStageRegFileWrite_payload_address[8]), .A2(n2616), 
        .B1(_zz_lastStageRegFileWrite_payload_address[9]), .B2(n2615), .ZN(
        n228) );
  aoi221d1 U793 ( .B1(n2615), .B2(_zz_lastStageRegFileWrite_payload_address[9]), .C1(n2616), .C2(_zz_lastStageRegFileWrite_payload_address[8]), .A(n228), 
        .ZN(n232) );
  oai22d1 U794 ( .A1(_zz_lastStageRegFileWrite_payload_address[11]), .A2(n2613), .B1(_zz_lastStageRegFileWrite_payload_address[10]), .B2(n2614), .ZN(n229) );
  aoi221d1 U795 ( .B1(n2614), .B2(
        _zz_lastStageRegFileWrite_payload_address[10]), .C1(n2613), .C2(
        _zz_lastStageRegFileWrite_payload_address[11]), .A(n229), .ZN(n231) );
  inv0d0 U796 ( .I(_zz_lastStageRegFileWrite_payload_address[7]), .ZN(n3316)
         );
  aoi22d1 U797 ( .A1(_zz_lastStageRegFileWrite_payload_address[7]), .A2(n2617), 
        .B1(\_zz__zz_decode_ENV_CTRL_2_1[20] ), .B2(n3316), .ZN(n230) );
  oai22d1 U798 ( .A1(n2613), .A2(
        HazardSimplePlugin_writeBackBuffer_payload_address[4]), .B1(n2616), 
        .B2(HazardSimplePlugin_writeBackBuffer_payload_address[1]), .ZN(n233)
         );
  aoi221d1 U799 ( .B1(n2613), .B2(
        HazardSimplePlugin_writeBackBuffer_payload_address[4]), .C1(
        HazardSimplePlugin_writeBackBuffer_payload_address[1]), .C2(n2616), 
        .A(n233), .ZN(n238) );
  inv0d0 U800 ( .I(HazardSimplePlugin_writeBackBuffer_payload_address[0]), 
        .ZN(n235) );
  oai22d1 U801 ( .A1(n2614), .A2(
        HazardSimplePlugin_writeBackBuffer_payload_address[3]), .B1(n235), 
        .B2(\_zz__zz_decode_ENV_CTRL_2_1[20] ), .ZN(n234) );
  aoi221d1 U802 ( .B1(n2614), .B2(
        HazardSimplePlugin_writeBackBuffer_payload_address[3]), .C1(
        \_zz__zz_decode_ENV_CTRL_2_1[20] ), .C2(n235), .A(n234), .ZN(n237) );
  aoim22d1 U803 ( .A1(HazardSimplePlugin_writeBackBuffer_payload_address[2]), 
        .A2(n2615), .B1(n2615), .B2(
        HazardSimplePlugin_writeBackBuffer_payload_address[2]), .Z(n236) );
  oai211d1 U804 ( .C1(n242), .C2(n241), .A(n240), .B(n239), .ZN(n280) );
  inv0d0 U805 ( .I(memory_INSTRUCTION[8]), .ZN(n6739) );
  nd02d0 U806 ( .A1(memory_arbitration_isValid), .A2(
        memory_REGFILE_WRITE_VALID), .ZN(n243) );
  aoi221d1 U807 ( .B1(decode_INSTRUCTION[16]), .B2(n6739), .C1(n2623), .C2(
        memory_INSTRUCTION[8]), .A(n243), .ZN(n255) );
  oai22d1 U808 ( .A1(memory_INSTRUCTION[9]), .A2(n2622), .B1(
        memory_INSTRUCTION[7]), .B2(n2624), .ZN(n244) );
  aoi221d1 U809 ( .B1(n174), .B2(memory_INSTRUCTION[7]), .C1(n2622), .C2(
        memory_INSTRUCTION[9]), .A(n244), .ZN(n254) );
  inv0d0 U810 ( .I(decode_INSTRUCTION[18]), .ZN(n2619) );
  oai22d1 U811 ( .A1(memory_INSTRUCTION[11]), .A2(n2618), .B1(n2619), .B2(
        memory_INSTRUCTION[10]), .ZN(n245) );
  aoi221d1 U812 ( .B1(n2618), .B2(memory_INSTRUCTION[11]), .C1(n173), .C2(
        memory_INSTRUCTION[10]), .A(n245), .ZN(n253) );
  inv0d0 U813 ( .I(_zz_lastStageRegFileWrite_payload_address[9]), .ZN(n3315)
         );
  oai22d1 U814 ( .A1(n2623), .A2(_zz_lastStageRegFileWrite_payload_address[8]), 
        .B1(n3315), .B2(decode_INSTRUCTION[17]), .ZN(n246) );
  aoi221d1 U815 ( .B1(n2623), .B2(_zz_lastStageRegFileWrite_payload_address[8]), .C1(decode_INSTRUCTION[17]), .C2(n3315), .A(n246), .ZN(n250) );
  oai222d1 U816 ( .A1(_zz_lastStageRegFileWrite_payload_address[7]), .A2(n2624), .B1(n3316), .B2(decode_INSTRUCTION[15]), .C1(
        _zz_lastStageRegFileWrite_payload_address[11]), .C2(n2618), .ZN(n247)
         );
  aoi211d1 U817 ( .C1(_zz_lastStageRegFileWrite_payload_address[11]), .C2(
        n2618), .A(n248), .B(n247), .ZN(n249) );
  oai211d1 U818 ( .C1(_zz_lastStageRegFileWrite_payload_address[10]), .C2(n173), .A(n250), .B(n249), .ZN(n251) );
  aoi21d1 U819 ( .B1(_zz_lastStageRegFileWrite_payload_address[10]), .B2(n173), 
        .A(n251), .ZN(n252) );
  aoi31d1 U820 ( .B1(n255), .B2(n254), .B3(n253), .A(n252), .ZN(n278) );
  oai22d1 U821 ( .A1(HazardSimplePlugin_writeBackBuffer_payload_address[0]), 
        .A2(n2624), .B1(n2618), .B2(
        HazardSimplePlugin_writeBackBuffer_payload_address[4]), .ZN(n256) );
  aoi221d1 U822 ( .B1(n174), .B2(
        HazardSimplePlugin_writeBackBuffer_payload_address[0]), .C1(n2618), 
        .C2(HazardSimplePlugin_writeBackBuffer_payload_address[4]), .A(n256), 
        .ZN(n260) );
  oai22d1 U823 ( .A1(HazardSimplePlugin_writeBackBuffer_payload_address[2]), 
        .A2(n2622), .B1(HazardSimplePlugin_writeBackBuffer_payload_address[3]), 
        .B2(n2619), .ZN(n257) );
  aoi221d1 U824 ( .B1(n173), .B2(
        HazardSimplePlugin_writeBackBuffer_payload_address[3]), .C1(n2622), 
        .C2(HazardSimplePlugin_writeBackBuffer_payload_address[2]), .A(n257), 
        .ZN(n259) );
  aoim22d1 U825 ( .A1(HazardSimplePlugin_writeBackBuffer_payload_address[1]), 
        .A2(n2623), .B1(n2623), .B2(
        HazardSimplePlugin_writeBackBuffer_payload_address[1]), .Z(n258) );
  nr02d0 U826 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[6]), .A2(
        _zz_decode_LEGAL_INSTRUCTION_1[2]), .ZN(n2555) );
  nr02d0 U827 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[4]), .A2(
        _zz_decode_LEGAL_INSTRUCTION_1[3]), .ZN(n2565) );
  aoi211d1 U828 ( .C1(n2585), .C2(n2578), .A(n2555), .B(n2565), .ZN(n276) );
  inv0d0 U829 ( .I(_zz__zz_execute_SRC2_3[1]), .ZN(n6738) );
  aoi22d1 U830 ( .A1(_zz__zz_execute_SRC2_3[1]), .A2(decode_INSTRUCTION_21), 
        .B1(n2616), .B2(n6738), .ZN(n272) );
  oai22d1 U831 ( .A1(_zz__zz_execute_SRC2_3[0]), .A2(n2617), .B1(
        _zz__zz_execute_SRC2_3[4]), .B2(n2613), .ZN(n261) );
  aoi221d1 U832 ( .B1(n2613), .B2(_zz__zz_execute_SRC2_3[4]), .C1(n2617), .C2(
        _zz__zz_execute_SRC2_3[0]), .A(n261), .ZN(n264) );
  aoi22d1 U833 ( .A1(_zz__zz_execute_SRC2_3[2]), .A2(n2615), .B1(
        decode_INSTRUCTION_22), .B2(n6722), .ZN(n263) );
  aoi22d1 U834 ( .A1(_zz__zz_execute_SRC2_3[3]), .A2(n2614), .B1(
        decode_INSTRUCTION_23), .B2(n6709), .ZN(n262) );
  oai22d1 U835 ( .A1(_zz__zz_execute_SRC2_3[4]), .A2(n2618), .B1(n2619), .B2(
        _zz__zz_execute_SRC2_3[3]), .ZN(n265) );
  aoi221d1 U836 ( .B1(n2618), .B2(_zz__zz_execute_SRC2_3[4]), .C1(n2619), .C2(
        _zz__zz_execute_SRC2_3[3]), .A(n265), .ZN(n269) );
  aoi22d1 U837 ( .A1(decode_INSTRUCTION[16]), .A2(n6738), .B1(
        _zz__zz_execute_SRC2_3[1]), .B2(n2623), .ZN(n268) );
  aoi22d1 U838 ( .A1(_zz__zz_execute_SRC2_3[2]), .A2(n2622), .B1(
        decode_INSTRUCTION[17]), .B2(n6722), .ZN(n267) );
  inv0d0 U839 ( .I(_zz__zz_execute_SRC2_3[0]), .ZN(n6753) );
  aoi22d1 U840 ( .A1(_zz__zz_execute_SRC2_3[0]), .A2(n2624), .B1(
        decode_INSTRUCTION[15]), .B2(n6753), .ZN(n266) );
  oai22d1 U841 ( .A1(n272), .A2(n271), .B1(n276), .B2(n270), .ZN(n274) );
  aoi31d1 U842 ( .B1(execute_arbitration_isValid), .B2(
        execute_REGFILE_WRITE_VALID), .B3(n274), .A(n273), .ZN(n275) );
  aon211d1 U843 ( .C1(n278), .C2(n277), .B(n276), .A(n275), .ZN(n279) );
  aon211d1 U844 ( .C1(n281), .C2(n280), .B(n279), .A(n2360), .ZN(n282) );
  nd04d1 U845 ( .A1(n2589), .A2(n284), .A3(n283), .A4(n282), .ZN(n2374) );
  inv0d0 U846 ( .I(n2374), .ZN(n3818) );
  inv0d0 U847 ( .I(n2474), .ZN(n2428) );
  nd02d0 U848 ( .A1(n2403), .A2(n2137), .ZN(n2214) );
  aoi211d1 U849 ( .C1(n2427), .C2(n2428), .A(n2198), .B(n2214), .ZN(n2050) );
  nr02d0 U850 ( .A1(reset), .A2(n2053), .ZN(n2358) );
  inv0d0 U851 ( .I(n2358), .ZN(n2355) );
  nr03d0 U852 ( .A1(n3818), .A2(n2054), .A3(n2355), .ZN(N1781) );
  buffd1 U853 ( .I(clk), .Z(n7254) );
  buffd1 U854 ( .I(n7254), .Z(n7208) );
  buffd1 U855 ( .I(n7208), .Z(n7206) );
  buffd1 U856 ( .I(n7208), .Z(n7234) );
  buffd1 U857 ( .I(n7234), .Z(n7235) );
  buffd1 U858 ( .I(n7123), .Z(n7211) );
  buffd1 U859 ( .I(n7235), .Z(n7210) );
  buffd1 U860 ( .I(n7210), .Z(n7212) );
  buffd1 U861 ( .I(n7235), .Z(n7209) );
  buffd1 U862 ( .I(n7123), .Z(n7207) );
  buffd1 U863 ( .I(n7234), .Z(n7205) );
  buffd1 U864 ( .I(clk), .Z(n7252) );
  buffd1 U865 ( .I(n7252), .Z(n7231) );
  buffd1 U866 ( .I(n7231), .Z(n7229) );
  buffd1 U867 ( .I(n7229), .Z(n7227) );
  buffd1 U868 ( .I(n7231), .Z(n7222) );
  buffd3 U869 ( .I(n7222), .Z(n7223) );
  buffd1 U870 ( .I(n7231), .Z(n7230) );
  buffd1 U871 ( .I(n7230), .Z(n7225) );
  buffd1 U872 ( .I(n7230), .Z(n7226) );
  buffd1 U873 ( .I(n7226), .Z(n7224) );
  buffd1 U874 ( .I(clk), .Z(n7253) );
  buffd1 U875 ( .I(n7253), .Z(n7217) );
  buffd1 U876 ( .I(n7217), .Z(n7216) );
  buffd1 U877 ( .I(n7217), .Z(n7232) );
  buffd1 U878 ( .I(n7232), .Z(n7233) );
  buffd1 U879 ( .I(n7233), .Z(n7221) );
  buffd1 U880 ( .I(n7221), .Z(n7219) );
  buffd1 U881 ( .I(n7232), .Z(n7213) );
  buffd1 U882 ( .I(n7217), .Z(n7214) );
  buffd1 U883 ( .I(n7221), .Z(n7215) );
  buffd1 U884 ( .I(n7233), .Z(n7218) );
  buffd1 U885 ( .I(n7218), .Z(n7220) );
  buffd1 U886 ( .I(clk), .Z(n7258) );
  buffd1 U887 ( .I(n7258), .Z(n7172) );
  buffd1 U888 ( .I(n7172), .Z(n7170) );
  buffd1 U889 ( .I(clk), .Z(n7260) );
  buffd1 U890 ( .I(n7260), .Z(n7154) );
  buffd1 U891 ( .I(n7154), .Z(n7246) );
  buffd1 U892 ( .I(n7246), .Z(n7151) );
  buffd1 U893 ( .I(n7154), .Z(n7152) );
  buffd1 U894 ( .I(n7246), .Z(n7247) );
  buffd1 U895 ( .I(n7247), .Z(n7155) );
  buffd1 U896 ( .I(n7247), .Z(n7159) );
  buffd1 U897 ( .I(n7159), .Z(n7157) );
  buffd1 U898 ( .I(n7159), .Z(n7153) );
  buffd1 U899 ( .I(clk), .Z(n7261) );
  buffd1 U900 ( .I(n7261), .Z(n7145) );
  buffd1 U901 ( .I(n7145), .Z(n7248) );
  buffd1 U902 ( .I(n7248), .Z(n7249) );
  buffd1 U903 ( .I(n7249), .Z(n7150) );
  buffd1 U904 ( .I(n7150), .Z(n7144) );
  buffd1 U905 ( .I(clk), .Z(n7259) );
  buffd1 U906 ( .I(n7259), .Z(n7163) );
  buffd1 U907 ( .I(n7163), .Z(n7244) );
  buffd1 U908 ( .I(n7244), .Z(n7245) );
  buffd1 U909 ( .I(n7245), .Z(n7164) );
  buffd1 U910 ( .I(n7150), .Z(n7148) );
  buffd1 U911 ( .I(n7249), .Z(n7146) );
  buffd1 U912 ( .I(n7247), .Z(n7156) );
  buffd1 U913 ( .I(n7156), .Z(n7158) );
  buffd1 U914 ( .I(n7145), .Z(n7143) );
  buffd1 U915 ( .I(n7248), .Z(n7142) );
  buffd1 U916 ( .I(n7244), .Z(n7160) );
  buffd1 U917 ( .I(n7245), .Z(n7168) );
  buffd1 U918 ( .I(n7168), .Z(n7166) );
  buffd1 U919 ( .I(n7245), .Z(n7165) );
  buffd1 U920 ( .I(n7165), .Z(n7167) );
  buffd1 U921 ( .I(n7249), .Z(n7147) );
  buffd1 U922 ( .I(n7147), .Z(n7149) );
  buffd1 U923 ( .I(n7163), .Z(n7161) );
  buffd1 U924 ( .I(n7168), .Z(n7162) );
  buffd1 U925 ( .I(n7231), .Z(n7228) );
  buffd1 U926 ( .I(clk), .Z(n7256) );
  buffd1 U927 ( .I(n7256), .Z(n7190) );
  buffd1 U928 ( .I(n7190), .Z(n7188) );
  buffd1 U929 ( .I(n7190), .Z(n7238) );
  buffd1 U930 ( .I(n7238), .Z(n7239) );
  buffd1 U931 ( .I(n7239), .Z(n7191) );
  buffd1 U932 ( .I(n7239), .Z(n7195) );
  buffd1 U933 ( .I(n7195), .Z(n7189) );
  buffd1 U934 ( .I(n7195), .Z(n7193) );
  buffd1 U935 ( .I(n7239), .Z(n7192) );
  buffd1 U936 ( .I(n7192), .Z(n7194) );
  buffd1 U937 ( .I(clk), .Z(n7255) );
  buffd1 U938 ( .I(n7255), .Z(n7199) );
  buffd1 U939 ( .I(n7199), .Z(n7236) );
  buffd1 U940 ( .I(n7236), .Z(n7237) );
  buffd1 U941 ( .I(n7237), .Z(n7204) );
  buffd1 U942 ( .I(n7204), .Z(n7198) );
  buffd1 U943 ( .I(n7204), .Z(n7202) );
  buffd1 U944 ( .I(n7237), .Z(n7201) );
  buffd1 U945 ( .I(n7201), .Z(n7203) );
  buffd1 U946 ( .I(n7236), .Z(n7196) );
  buffd1 U947 ( .I(n7199), .Z(n7197) );
  buffd1 U948 ( .I(n7237), .Z(n7200) );
  buffd1 U949 ( .I(clk), .Z(n7262) );
  buffd1 U950 ( .I(n7262), .Z(n7136) );
  buffd1 U951 ( .I(n7136), .Z(n7250) );
  buffd1 U952 ( .I(n7250), .Z(n7251) );
  buffd1 U953 ( .I(n7251), .Z(n7137) );
  buffd1 U954 ( .I(n7172), .Z(n7242) );
  buffd1 U955 ( .I(n7242), .Z(n7169) );
  buffd1 U956 ( .I(clk), .Z(n7263) );
  buffd3 U957 ( .I(n7263), .Z(n7123) );
  buffd1 U958 ( .I(n7123), .Z(n7125) );
  buffd1 U959 ( .I(n7125), .Z(n7130) );
  buffd1 U960 ( .I(n7123), .Z(n7124) );
  buffd1 U961 ( .I(n7124), .Z(n7128) );
  buffd1 U962 ( .I(n7128), .Z(n7132) );
  buffd1 U963 ( .I(n7242), .Z(n7243) );
  buffd1 U964 ( .I(n7243), .Z(n7174) );
  buffd1 U965 ( .I(n7174), .Z(n7176) );
  buffd1 U966 ( .I(n7128), .Z(n7127) );
  buffd1 U967 ( .I(n7123), .Z(n7129) );
  buffd1 U968 ( .I(n7243), .Z(n7177) );
  buffd1 U969 ( .I(n7177), .Z(n7175) );
  buffd1 U970 ( .I(n7177), .Z(n7171) );
  buffd1 U971 ( .I(n7243), .Z(n7173) );
  buffd1 U972 ( .I(n7263), .Z(n7131) );
  buffd1 U973 ( .I(n7124), .Z(n7126) );
  buffd1 U974 ( .I(n7251), .Z(n7138) );
  buffd1 U975 ( .I(n7138), .Z(n7140) );
  buffd1 U976 ( .I(n7251), .Z(n7141) );
  buffd1 U977 ( .I(n7141), .Z(n7135) );
  buffd1 U978 ( .I(clk), .Z(n7257) );
  buffd1 U979 ( .I(n7257), .Z(n7181) );
  buffd1 U980 ( .I(n7181), .Z(n7240) );
  buffd1 U981 ( .I(n7240), .Z(n7241) );
  buffd1 U982 ( .I(n7241), .Z(n7186) );
  buffd1 U983 ( .I(n7186), .Z(n7184) );
  buffd1 U984 ( .I(n7241), .Z(n7183) );
  buffd1 U985 ( .I(n7183), .Z(n7185) );
  buffd1 U986 ( .I(n7141), .Z(n7139) );
  buffd1 U987 ( .I(n7240), .Z(n7178) );
  buffd1 U988 ( .I(n7241), .Z(n7182) );
  buffd1 U989 ( .I(n7181), .Z(n7179) );
  buffd1 U990 ( .I(n7250), .Z(n7133) );
  buffd1 U991 ( .I(n7136), .Z(n7134) );
  buffd1 U992 ( .I(n7238), .Z(n7187) );
  buffd1 U993 ( .I(n7186), .Z(n7180) );
  buffd1 U994 ( .I(n3235), .Z(n3232) );
  buffd1 U995 ( .I(n3232), .Z(n3247) );
  buffd1 U996 ( .I(n3247), .Z(n3238) );
  aoim22d1 U997 ( .A1(n6738), .A2(n3235), .B1(n3238), .B2(decode_INSTRUCTION_8), .Z(n5954) );
  nr02d0 U998 ( .A1(dBus_cmd_halfPipe_payload_address[1]), .A2(
        dBus_cmd_halfPipe_payload_address[0]), .ZN(n366) );
  nd12d0 U999 ( .A1(n366), .A2(dBusWishbone_WE), .ZN(dBusWishbone_SEL[0]) );
  nr03d0 U1000 ( .A1(dBus_cmd_halfPipe_payload_address[0]), .A2(
        dBus_cmd_halfPipe_payload_size[0]), .A3(
        dBus_cmd_halfPipe_payload_size[1]), .ZN(n367) );
  oai21d1 U1001 ( .B1(dBus_cmd_halfPipe_payload_address[1]), .B2(n367), .A(
        dBusWishbone_WE), .ZN(dBusWishbone_SEL[1]) );
  an02d0 U1002 ( .A1(_zz_CsrPlugin_csrMapping_readDataInit[7]), .A2(
        externalInterruptArray_regNext[7]), .Z(n2307) );
  nd02d0 U1003 ( .A1(_zz_CsrPlugin_csrMapping_readDataInit[3]), .A2(
        externalInterruptArray_regNext[3]), .ZN(n288) );
  nd02d0 U1004 ( .A1(_zz_CsrPlugin_csrMapping_readDataInit[2]), .A2(
        externalInterruptArray_regNext[2]), .ZN(n287) );
  nd02d0 U1005 ( .A1(_zz_CsrPlugin_csrMapping_readDataInit[0]), .A2(
        externalInterruptArray_regNext[0]), .ZN(n2247) );
  nd02d0 U1006 ( .A1(_zz_CsrPlugin_csrMapping_readDataInit[1]), .A2(
        externalInterruptArray_regNext[1]), .ZN(n286) );
  aoi211d1 U1007 ( .C1(_zz_CsrPlugin_csrMapping_readDataInit[6]), .C2(
        externalInterruptArray_regNext[6]), .A(n2307), .B(n289), .ZN(n292) );
  nd02d0 U1008 ( .A1(_zz_CsrPlugin_csrMapping_readDataInit[4]), .A2(
        externalInterruptArray_regNext[4]), .ZN(n291) );
  nd02d0 U1009 ( .A1(_zz_CsrPlugin_csrMapping_readDataInit[5]), .A2(
        externalInterruptArray_regNext[5]), .ZN(n290) );
  nr02d0 U1010 ( .A1(\IBusCachedPlugin_cache/_zz_ways_0_tags_port[0] ), .A2(
        \IBusCachedPlugin_cache/lineLoader_flushCounter[0] ), .ZN(n3060) );
  inv0d0 U1011 ( .I(_zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1), 
        .ZN(n2372) );
  nd03d0 U1012 ( .A1(\IBusCachedPlugin_cache/lineLoader_flushPending ), .A2(
        n2372), .A3(n2413), .ZN(n2410) );
  inv0d0 U1013 ( .I(n2410), .ZN(n293) );
  nd02d0 U1014 ( .A1(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[1] ), 
        .A2(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[2] ), 
        .ZN(n3138) );
  nd02d0 U1015 ( .A1(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[0] ), 
        .A2(iBus_rsp_valid), .ZN(n2407) );
  nr02d0 U1016 ( .A1(n3138), .A2(n2407), .ZN(n2414) );
  aoi21d1 U1017 ( .B1(iBusWishbone_ACK), .B2(
        \IBusCachedPlugin_cache/lineLoader_valid ), .A(
        \IBusCachedPlugin_cache/lineLoader_cmdSent ), .ZN(n294) );
  nr03d0 U1018 ( .A1(n2412), .A2(n2414), .A3(n294), .ZN(n6082) );
  nd02d0 U1019 ( .A1(iBusWishbone_ACK), .A2(when_InstructionCache_l239), .ZN(
        n2219) );
  inv0d0 U1020 ( .I(n7113), .ZN(n6740) );
  inv0d0 U1021 ( .I(execute_INSTRUCTION[5]), .ZN(n6781) );
  inv0d0 U1022 ( .I(n561), .ZN(n2335) );
  aoi22d1 U1023 ( .A1(n6740), .A2(CsrPlugin_pipelineLiberator_pcValids_1), 
        .B1(CsrPlugin_pipelineLiberator_pcValids_0), .B2(n6996), .ZN(n296) );
  nr02d0 U1024 ( .A1(n2335), .A2(n296), .ZN(n6132) );
  inv0d0 U1025 ( .I(n299), .ZN(n2942) );
  or02d0 U1026 ( .A1(n299), .A2(n562), .Z(n2748) );
  inv0d1 U1027 ( .I(n2748), .ZN(n2872) );
  inv0d0 U1028 ( .I(execute_CsrPlugin_csr_835), .ZN(n2538) );
  inv0d1 U1029 ( .I(n2538), .ZN(n2327) );
  aoi22d1 U1030 ( .A1(execute_CsrPlugin_csr_3008), .A2(
        _zz_CsrPlugin_csrMapping_readDataInit[12]), .B1(n2327), .B2(
        CsrPlugin_mtval[12]), .ZN(n298) );
  aoi22d1 U1031 ( .A1(CsrPlugin_mepc[12]), .A2(execute_CsrPlugin_csr_833), 
        .B1(execute_CsrPlugin_csr_768), .B2(CsrPlugin_mstatus_MPP[1]), .ZN(
        n297) );
  nd02d0 U1032 ( .A1(n298), .A2(n297), .ZN(n2294) );
  inv0d0 U1033 ( .I(n299), .ZN(n2749) );
  aoi22d1 U1034 ( .A1(n2872), .A2(n2294), .B1(memory_REGFILE_WRITE_DATA[12]), 
        .B2(n3020), .ZN(n325) );
  inv0d0 U1035 ( .I(n300), .ZN(n2640) );
  nr03d1 U1036 ( .A1(execute_LightShifterPlugin_isActive), .A2(
        execute_SHIFT_CTRL[1]), .A3(n2640), .ZN(n2969) );
  inv0d0 U1037 ( .I(execute_RS1[11]), .ZN(n6285) );
  nr02d0 U1038 ( .A1(n2111), .A2(n6285), .ZN(n2873) );
  inv0d0 U1039 ( .I(execute_ALU_CTRL[0]), .ZN(n2588) );
  nd02d0 U1040 ( .A1(execute_ALU_CTRL[1]), .A2(n2588), .ZN(n301) );
  oai211d1 U1041 ( .C1(execute_ALU_CTRL[1]), .C2(n2588), .A(n2640), .B(n301), 
        .ZN(n3005) );
  inv0d0 U1042 ( .I(execute_RS1[12]), .ZN(n6282) );
  oai22d1 U1043 ( .A1(n336), .A2(n6282), .B1(n6681), .B2(n302), .ZN(n2869) );
  aoi22d1 U1044 ( .A1(n2109), .A2(execute_RS2[12]), .B1(n2105), .B2(
        execute_PC[12]), .ZN(n306) );
  buffd1 U1045 ( .I(_zz__zz_execute_SRC2_3[11]), .Z(n6343) );
  nd02d0 U1046 ( .A1(n306), .A2(n305), .ZN(n319) );
  aoim22d1 U1047 ( .A1(execute_SRC_USE_SUB_LESS), .A2(n319), .B1(n319), .B2(
        execute_SRC_USE_SUB_LESS), .Z(n340) );
  aoi22d1 U1048 ( .A1(n2109), .A2(execute_RS2[11]), .B1(n2105), .B2(
        execute_PC[11]), .ZN(n307) );
  nd02d0 U1049 ( .A1(n307), .A2(n305), .ZN(n2874) );
  aoim22d1 U1050 ( .A1(execute_SRC_USE_SUB_LESS), .A2(n2874), .B1(n2874), .B2(
        n2117), .Z(n2865) );
  inv0d0 U1051 ( .I(execute_RS1[10]), .ZN(n6286) );
  nr02d0 U1052 ( .A1(n2111), .A2(n6286), .ZN(n2885) );
  aoi222d1 U1053 ( .A1(n308), .A2(_zz__zz_execute_SRC2_3[10]), .B1(n2105), 
        .B2(execute_PC[10]), .C1(n2114), .C2(execute_RS2[10]), .ZN(n2890) );
  aoim22d1 U1054 ( .A1(n2890), .A2(n2594), .B1(n2110), .B2(n2890), .Z(n2883)
         );
  inv0d0 U1055 ( .I(execute_RS1[9]), .ZN(n6287) );
  nr02d0 U1056 ( .A1(n2111), .A2(n6287), .ZN(n2899) );
  aoi222d1 U1057 ( .A1(n308), .A2(_zz__zz_execute_SRC2_3[9]), .B1(n2105), .B2(
        execute_PC[9]), .C1(n2114), .C2(execute_RS2[9]), .ZN(n2906) );
  aoim22d1 U1058 ( .A1(n2906), .A2(n2594), .B1(n2110), .B2(n2906), .Z(n2896)
         );
  inv0d0 U1059 ( .I(execute_RS1[8]), .ZN(n6288) );
  nr02d0 U1060 ( .A1(n2111), .A2(n6288), .ZN(n2914) );
  aoi222d1 U1061 ( .A1(n308), .A2(_zz__zz_execute_SRC2_3[8]), .B1(n2113), .B2(
        execute_PC[8]), .C1(n2114), .C2(execute_RS2[8]), .ZN(n2920) );
  aoim22d1 U1062 ( .A1(n2920), .A2(n2594), .B1(n2110), .B2(n2920), .Z(n2912)
         );
  inv0d0 U1063 ( .I(execute_RS1[7]), .ZN(n6289) );
  nr02d0 U1064 ( .A1(n336), .A2(n6289), .ZN(n2931) );
  aoi222d1 U1065 ( .A1(n308), .A2(_zz__zz_execute_SRC2_3[7]), .B1(n2105), .B2(
        execute_PC[7]), .C1(n2114), .C2(execute_RS2[7]), .ZN(n2934) );
  aoim22d1 U1066 ( .A1(n2934), .A2(n2594), .B1(n2110), .B2(n2934), .Z(n2929)
         );
  inv0d0 U1067 ( .I(execute_RS1[6]), .ZN(n6291) );
  aoi222d1 U1068 ( .A1(n308), .A2(_zz__zz_execute_SRC2_3[6]), .B1(n2105), .B2(
        execute_PC[6]), .C1(n2114), .C2(execute_RS2[6]), .ZN(n2947) );
  aoim22d1 U1069 ( .A1(n2947), .A2(n2594), .B1(n2110), .B2(n2947), .Z(n2949)
         );
  inv0d0 U1070 ( .I(execute_RS1[5]), .ZN(n6292) );
  nr02d0 U1071 ( .A1(n336), .A2(n6292), .ZN(n2965) );
  aoi222d1 U1072 ( .A1(n308), .A2(_zz__zz_execute_SRC2_3[5]), .B1(n2113), .B2(
        execute_PC[5]), .C1(n2114), .C2(execute_RS2[5]), .ZN(n2975) );
  aoim22d1 U1073 ( .A1(n2975), .A2(n2594), .B1(n2110), .B2(n2975), .Z(n2963)
         );
  inv0d0 U1074 ( .I(execute_RS1[4]), .ZN(n6294) );
  inv0d0 U1075 ( .I(_zz__zz_execute_SRC1_1[4]), .ZN(n6269) );
  oai22d1 U1076 ( .A1(n336), .A2(n6294), .B1(n309), .B2(n6269), .ZN(n2990) );
  inv0d0 U1077 ( .I(n2988), .ZN(n2986) );
  aoi22d1 U1078 ( .A1(n2986), .A2(n2110), .B1(n2117), .B2(n2988), .ZN(n2977)
         );
  inv0d0 U1079 ( .I(execute_RS1[3]), .ZN(n6296) );
  inv0d0 U1080 ( .I(_zz__zz_execute_SRC1_1[3]), .ZN(n6271) );
  oai22d1 U1081 ( .A1(n2111), .A2(n6296), .B1(n309), .B2(n6271), .ZN(n563) );
  aoi22d1 U1082 ( .A1(n353), .A2(n2110), .B1(n2117), .B2(n361), .ZN(n355) );
  inv0d0 U1083 ( .I(execute_RS1[2]), .ZN(n6300) );
  nr02d0 U1084 ( .A1(_zz__zz_execute_SRC1_1[2]), .A2(n2597), .ZN(n332) );
  oan211d1 U1085 ( .C1(execute_SRC1_CTRL[0]), .C2(n6300), .B(n2601), .A(n332), 
        .ZN(n3016) );
  inv0d0 U1086 ( .I(n3000), .ZN(n3015) );
  aoi22d1 U1087 ( .A1(n3000), .A2(n2110), .B1(n2117), .B2(n3015), .ZN(n3002)
         );
  aoi22d1 U1088 ( .A1(n2932), .A2(n2869), .B1(n312), .B2(n3003), .ZN(n6897) );
  nr02d0 U1089 ( .A1(n2572), .A2(n315), .ZN(n313) );
  inv0d1 U1090 ( .I(n314), .ZN(n2870) );
  inv0d0 U1091 ( .I(execute_RS1[13]), .ZN(n6280) );
  oai22d1 U1092 ( .A1(n336), .A2(n6280), .B1(n6666), .B2(n302), .ZN(n2291) );
  nr03d0 U1093 ( .A1(n3679), .A2(n2572), .A3(n315), .ZN(n2818) );
  inv0d0 U1094 ( .I(n2818), .ZN(n2980) );
  inv0d1 U1095 ( .I(n2980), .ZN(n3027) );
  aoi22d1 U1096 ( .A1(n2870), .A2(n2291), .B1(n3027), .B2(
        memory_REGFILE_WRITE_DATA[13]), .ZN(n317) );
  nd03d0 U1097 ( .A1(execute_ALU_CTRL[1]), .A2(n2640), .A3(n2588), .ZN(n320)
         );
  nd13d1 U1098 ( .A1(n320), .A2(execute_ALU_BITWISE_CTRL[0]), .A3(n6681), .ZN(
        n3006) );
  inv0d2 U1099 ( .I(n3006), .ZN(n3026) );
  nr03d0 U1100 ( .A1(execute_SHIFT_CTRL[1]), .A2(n3679), .A3(n2640), .ZN(n2984) );
  inv0d0 U1101 ( .I(n2984), .ZN(n2943) );
  inv0d1 U1102 ( .I(n2943), .ZN(n3029) );
  aoi22d1 U1103 ( .A1(n3026), .A2(n319), .B1(n3029), .B2(
        memory_REGFILE_WRITE_DATA[11]), .ZN(n316) );
  oai211d1 U1104 ( .C1(n3005), .C2(n6897), .A(n317), .B(n316), .ZN(n318) );
  inv0d0 U1105 ( .I(n3033), .ZN(n2856) );
  aon211d1 U1106 ( .C1(n2969), .C2(n2873), .B(n318), .A(n2856), .ZN(n324) );
  nr03d0 U1107 ( .A1(n320), .A2(n6681), .A3(execute_ALU_BITWISE_CTRL[0]), .ZN(
        n2761) );
  inv0d0 U1108 ( .I(n2761), .ZN(n2961) );
  nr02d1 U1109 ( .A1(n2996), .A2(n2961), .ZN(n3040) );
  nr02d1 U1110 ( .A1(n2996), .A2(n3006), .ZN(n2989) );
  aon211d1 U1111 ( .C1(n3040), .C2(n319), .B(n2989), .A(n2869), .ZN(n323) );
  inv0d0 U1112 ( .I(n2869), .ZN(n2293) );
  mx02d1 U1113 ( .I0(n2869), .I1(n2293), .S(n319), .Z(n3756) );
  nr02d0 U1114 ( .A1(execute_ALU_BITWISE_CTRL[0]), .A2(n6681), .ZN(n321) );
  aoi211d1 U1115 ( .C1(execute_ALU_BITWISE_CTRL[0]), .C2(n6681), .A(n321), .B(
        n320), .ZN(n2960) );
  buffd1 U1116 ( .I(n2960), .Z(n3032) );
  inv0d0 U1117 ( .I(n3032), .ZN(n3013) );
  nr02d1 U1118 ( .A1(n2996), .A2(n3013), .ZN(n2994) );
  nd02d0 U1119 ( .A1(n3756), .A2(n2994), .ZN(n322) );
  inv0d0 U1120 ( .I(execute_RS1[22]), .ZN(n6265) );
  inv0d0 U1121 ( .I(_zz__zz_execute_BranchPlugin_branch_src2_1), .ZN(n6298) );
  oai22d1 U1122 ( .A1(n336), .A2(n6265), .B1(n6298), .B2(n302), .ZN(n2775) );
  inv0d0 U1123 ( .I(n2775), .ZN(n2752) );
  aoi22d1 U1124 ( .A1(n2109), .A2(execute_RS2[22]), .B1(n2113), .B2(
        execute_PC[22]), .ZN(n326) );
  nd02d0 U1125 ( .A1(n326), .A2(n305), .ZN(n345) );
  mx02d1 U1126 ( .I0(n2775), .I1(n2752), .S(n345), .Z(n3757) );
  inv0d0 U1127 ( .I(memory_REGFILE_WRITE_DATA[22]), .ZN(n2764) );
  inv0d0 U1128 ( .I(execute_CsrPlugin_csr_3008), .ZN(n2244) );
  inv0d1 U1129 ( .I(n2244), .ZN(n2328) );
  aoi222d1 U1130 ( .A1(CsrPlugin_mepc[22]), .A2(execute_CsrPlugin_csr_833), 
        .B1(n2328), .B2(_zz_CsrPlugin_csrMapping_readDataInit[22]), .C1(n2327), 
        .C2(CsrPlugin_mtval[22]), .ZN(n2268) );
  oai22d1 U1131 ( .A1(n2749), .A2(n2764), .B1(n2268), .B2(n2748), .ZN(n327) );
  aoi21d1 U1132 ( .B1(n3757), .B2(n2994), .A(n327), .ZN(n348) );
  inv0d0 U1133 ( .I(execute_RS1[21]), .ZN(n6266) );
  inv0d0 U1134 ( .I(_zz__zz_execute_BranchPlugin_branch_src2_0), .ZN(n6303) );
  oai22d1 U1135 ( .A1(n336), .A2(n6266), .B1(n6303), .B2(n302), .ZN(n2782) );
  aoim22d1 U1136 ( .A1(execute_SRC_USE_SUB_LESS), .A2(n345), .B1(n345), .B2(
        n2117), .Z(n2119) );
  aoi22d1 U1137 ( .A1(n2114), .A2(execute_RS2[21]), .B1(n2113), .B2(
        execute_PC[21]), .ZN(n328) );
  nd02d0 U1138 ( .A1(n328), .A2(n305), .ZN(n2781) );
  inv0d0 U1139 ( .I(n2781), .ZN(n2774) );
  aoi22d1 U1140 ( .A1(n2774), .A2(n2110), .B1(n2117), .B2(n2781), .ZN(n2772)
         );
  inv0d0 U1141 ( .I(execute_RS1[20]), .ZN(n6267) );
  inv0d0 U1142 ( .I(_zz__zz_execute_BranchPlugin_branch_src2[10]), .ZN(n6307)
         );
  oai22d1 U1143 ( .A1(n2111), .A2(n6267), .B1(n6307), .B2(n302), .ZN(n2805) );
  aoi22d1 U1144 ( .A1(n2109), .A2(execute_RS2[20]), .B1(n2113), .B2(
        execute_PC[20]), .ZN(n329) );
  nd02d0 U1145 ( .A1(n329), .A2(n305), .ZN(n2797) );
  inv0d0 U1146 ( .I(n2797), .ZN(n2792) );
  aoi22d1 U1147 ( .A1(n2792), .A2(n2110), .B1(n2117), .B2(n2797), .ZN(n2788)
         );
  inv0d0 U1148 ( .I(execute_RS1[19]), .ZN(n6270) );
  oai22d1 U1149 ( .A1(n2111), .A2(n6270), .B1(n302), .B2(n6269), .ZN(n2812) );
  aoi22d1 U1150 ( .A1(n2114), .A2(execute_RS2[19]), .B1(n2113), .B2(
        execute_PC[19]), .ZN(n330) );
  nd02d0 U1151 ( .A1(n330), .A2(n305), .ZN(n2811) );
  aoim22d1 U1152 ( .A1(execute_SRC_USE_SUB_LESS), .A2(n2811), .B1(n2811), .B2(
        n2117), .Z(n2802) );
  inv0d0 U1153 ( .I(execute_RS1[18]), .ZN(n6272) );
  oai22d1 U1154 ( .A1(n2111), .A2(n6272), .B1(n302), .B2(n6271), .ZN(n2835) );
  aoi22d1 U1155 ( .A1(n2109), .A2(execute_RS2[18]), .B1(n2113), .B2(
        execute_PC[18]), .ZN(n331) );
  nd02d0 U1156 ( .A1(n331), .A2(n305), .ZN(n2824) );
  aoim22d1 U1157 ( .A1(execute_SRC_USE_SUB_LESS), .A2(n2824), .B1(n2824), .B2(
        n2117), .Z(n2816) );
  inv0d0 U1158 ( .I(execute_RS1[17]), .ZN(n6274) );
  aoi211d1 U1159 ( .C1(n2597), .C2(n6274), .A(execute_SRC1_CTRL[1]), .B(n332), 
        .ZN(n2838) );
  aoi22d1 U1160 ( .A1(n2109), .A2(execute_RS2[17]), .B1(n2105), .B2(
        execute_PC[17]), .ZN(n333) );
  nd02d0 U1161 ( .A1(n333), .A2(n305), .ZN(n2839) );
  aoim22d1 U1162 ( .A1(execute_SRC_USE_SUB_LESS), .A2(n2839), .B1(n2839), .B2(
        n2117), .Z(n2831) );
  inv0d0 U1163 ( .I(execute_RS1[16]), .ZN(n6276) );
  oai22d1 U1164 ( .A1(n2111), .A2(n6276), .B1(n6275), .B2(n302), .ZN(n2282) );
  aoi22d1 U1165 ( .A1(n2109), .A2(execute_RS2[16]), .B1(n2105), .B2(
        execute_PC[16]), .ZN(n334) );
  nd02d0 U1166 ( .A1(n334), .A2(n305), .ZN(n388) );
  aoim22d1 U1167 ( .A1(execute_SRC_USE_SUB_LESS), .A2(n388), .B1(n388), .B2(
        n2117), .Z(n383) );
  inv0d0 U1168 ( .I(execute_RS1[15]), .ZN(n6278) );
  oai22d1 U1169 ( .A1(n2111), .A2(n6278), .B1(n6277), .B2(n302), .ZN(n2848) );
  aoi22d1 U1170 ( .A1(n2109), .A2(execute_RS2[15]), .B1(n2113), .B2(
        execute_PC[15]), .ZN(n335) );
  nd02d0 U1171 ( .A1(n335), .A2(n305), .ZN(n400) );
  aoim22d1 U1172 ( .A1(execute_SRC_USE_SUB_LESS), .A2(n400), .B1(n400), .B2(
        n2117), .Z(n395) );
  inv0d0 U1173 ( .I(execute_RS1[14]), .ZN(n6279) );
  inv0d0 U1174 ( .I(_zz__zz_execute_BranchPlugin_branch_src2[13]), .ZN(n6650)
         );
  oai22d1 U1175 ( .A1(n336), .A2(n6279), .B1(n302), .B2(n6650), .ZN(n2863) );
  aoi22d1 U1176 ( .A1(n2109), .A2(execute_RS2[14]), .B1(n2113), .B2(
        execute_PC[14]), .ZN(n337) );
  nd02d0 U1177 ( .A1(n337), .A2(n305), .ZN(n2862) );
  aoim22d1 U1178 ( .A1(execute_SRC_USE_SUB_LESS), .A2(n2862), .B1(n2862), .B2(
        execute_SRC_USE_SUB_LESS), .Z(n2850) );
  aoi22d1 U1179 ( .A1(n2109), .A2(execute_RS2[13]), .B1(n2113), .B2(
        execute_PC[13]), .ZN(n338) );
  nd02d0 U1180 ( .A1(n338), .A2(n305), .ZN(n375) );
  aoim22d1 U1181 ( .A1(execute_SRC_USE_SUB_LESS), .A2(n375), .B1(n375), .B2(
        execute_SRC_USE_SUB_LESS), .Z(n370) );
  aoi22d1 U1182 ( .A1(n2932), .A2(n2775), .B1(n341), .B2(n2897), .ZN(n6846) );
  inv0d0 U1183 ( .I(execute_RS1[23]), .ZN(n6264) );
  inv0d0 U1184 ( .I(_zz__zz_execute_BranchPlugin_branch_src2_2), .ZN(n6295) );
  oai22d1 U1185 ( .A1(n2111), .A2(n6264), .B1(n6295), .B2(n302), .ZN(n2760) );
  aoi22d1 U1186 ( .A1(n2870), .A2(n2760), .B1(n3027), .B2(
        memory_REGFILE_WRITE_DATA[23]), .ZN(n343) );
  aoi22d1 U1187 ( .A1(n3026), .A2(n345), .B1(n3029), .B2(
        memory_REGFILE_WRITE_DATA[21]), .ZN(n342) );
  oai211d1 U1188 ( .C1(n3005), .C2(n6846), .A(n343), .B(n342), .ZN(n344) );
  aon211d1 U1189 ( .C1(n2969), .C2(n2782), .B(n344), .A(n2856), .ZN(n347) );
  aon211d1 U1190 ( .C1(n3040), .C2(n345), .B(n2989), .A(n2775), .ZN(n346) );
  inv0d1 U1191 ( .I(n2748), .ZN(n2999) );
  aoi22d1 U1192 ( .A1(n2327), .A2(CsrPlugin_mtval[3]), .B1(
        execute_CsrPlugin_csr_772), .B2(CsrPlugin_mie_MSIE), .ZN(n352) );
  aoi22d1 U1193 ( .A1(CsrPlugin_mepc[3]), .A2(execute_CsrPlugin_csr_833), .B1(
        execute_CsrPlugin_csr_834), .B2(CsrPlugin_mcause_exceptionCode[3]), 
        .ZN(n351) );
  aoi22d1 U1194 ( .A1(execute_CsrPlugin_csr_768), .A2(CsrPlugin_mstatus_MIE), 
        .B1(execute_CsrPlugin_csr_836), .B2(CsrPlugin_mip_MSIP), .ZN(n350) );
  aon211d1 U1195 ( .C1(execute_CsrPlugin_csr_4032), .C2(
        externalInterruptArray_regNext[3]), .B(execute_CsrPlugin_csr_3008), 
        .A(_zz_CsrPlugin_csrMapping_readDataInit[3]), .ZN(n349) );
  aoi22d1 U1196 ( .A1(n2999), .A2(n564), .B1(memory_REGFILE_WRITE_DATA[3]), 
        .B2(n3020), .ZN(n364) );
  inv0d0 U1197 ( .I(n563), .ZN(n3008) );
  aoi22d1 U1198 ( .A1(n353), .A2(n3008), .B1(n563), .B2(n361), .ZN(n3741) );
  inv0d0 U1199 ( .I(n3016), .ZN(n3023) );
  aoi22d1 U1200 ( .A1(n3026), .A2(n563), .B1(n2818), .B2(
        memory_REGFILE_WRITE_DATA[4]), .ZN(n359) );
  inv0d0 U1201 ( .I(n2990), .ZN(n2985) );
  aoi22d1 U1202 ( .A1(execute_SRC2_FORCE_ZERO), .A2(n563), .B1(n356), .B2(
        n3003), .ZN(n6964) );
  oai22d1 U1203 ( .A1(n2985), .A2(n314), .B1(n3005), .B2(n6964), .ZN(n357) );
  aoi21d1 U1204 ( .B1(n3029), .B2(memory_REGFILE_WRITE_DATA[2]), .A(n357), 
        .ZN(n358) );
  oai211d1 U1205 ( .C1(n3035), .C2(n3023), .A(n359), .B(n358), .ZN(n360) );
  aon211d1 U1206 ( .C1(n3032), .C2(n3741), .B(n360), .A(n2856), .ZN(n363) );
  aon211d1 U1207 ( .C1(n3040), .C2(n563), .B(n2989), .A(n361), .ZN(n362) );
  inv0d0 U1208 ( .I(dBus_cmd_halfPipe_payload_size[1]), .ZN(n6665) );
  inv0d0 U1209 ( .I(dBus_cmd_halfPipe_payload_address[1]), .ZN(n6982) );
  inv0d0 U1210 ( .I(dBus_cmd_halfPipe_payload_address[0]), .ZN(n6995) );
  oan211d1 U1211 ( .C1(dBus_cmd_halfPipe_payload_size[0]), .C2(
        dBus_cmd_halfPipe_payload_size[1]), .B(n6982), .A(n6995), .ZN(n365) );
  aon211d1 U1212 ( .C1(n366), .C2(n6665), .B(n365), .A(dBusWishbone_WE), .ZN(
        dBusWishbone_SEL[2]) );
  oai211d1 U1213 ( .C1(n367), .C2(n6982), .A(dBusWishbone_WE), .B(n6665), .ZN(
        dBusWishbone_SEL[3]) );
  inv0d0 U1214 ( .I(CsrPlugin_mepc[13]), .ZN(n3605) );
  aoi22d1 U1215 ( .A1(n2328), .A2(_zz_CsrPlugin_csrMapping_readDataInit[13]), 
        .B1(execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[13]), .ZN(n368) );
  oai21d1 U1216 ( .B1(n3605), .B2(n2541), .A(n368), .ZN(n2290) );
  aoi22d1 U1217 ( .A1(n2872), .A2(n2290), .B1(memory_REGFILE_WRITE_DATA[13]), 
        .B2(n3020), .ZN(n379) );
  inv0d0 U1218 ( .I(n2291), .ZN(n2855) );
  mx02d1 U1219 ( .I0(n2291), .I1(n2855), .S(n375), .Z(n3753) );
  aoi22d1 U1220 ( .A1(n2994), .A2(n3753), .B1(n2923), .B2(n2869), .ZN(n378) );
  inv0d0 U1221 ( .I(memory_REGFILE_WRITE_DATA[12]), .ZN(n2867) );
  inv0d0 U1222 ( .I(n2863), .ZN(n2860) );
  aoi22d1 U1223 ( .A1(n2932), .A2(n2291), .B1(n371), .B2(n3003), .ZN(n6896) );
  oai22d1 U1224 ( .A1(n2860), .A2(n314), .B1(n3005), .B2(n6896), .ZN(n372) );
  aoi31d1 U1225 ( .B1(n2761), .B2(n2291), .B3(n375), .A(n372), .ZN(n373) );
  oai21d1 U1226 ( .B1(n2943), .B2(n2867), .A(n373), .ZN(n374) );
  aon211d1 U1227 ( .C1(n3027), .C2(memory_REGFILE_WRITE_DATA[14]), .B(n374), 
        .A(n2856), .ZN(n377) );
  oai21d1 U1228 ( .B1(n2291), .B2(n375), .A(n2989), .ZN(n376) );
  inv0d0 U1229 ( .I(n2282), .ZN(n2842) );
  mx02d1 U1230 ( .I0(n2842), .I1(n2282), .S(n388), .Z(n3746) );
  inv0d0 U1231 ( .I(n3746), .ZN(n380) );
  aoi22d1 U1232 ( .A1(n2994), .A2(n380), .B1(n2923), .B2(n2848), .ZN(n392) );
  inv0d0 U1233 ( .I(CsrPlugin_mepc[16]), .ZN(n3614) );
  aoi22d1 U1234 ( .A1(n2328), .A2(_zz_CsrPlugin_csrMapping_readDataInit[16]), 
        .B1(n2327), .B2(CsrPlugin_mtval[16]), .ZN(n381) );
  oai21d1 U1235 ( .B1(n3614), .B2(n2541), .A(n381), .ZN(n2281) );
  aoi22d1 U1236 ( .A1(n2872), .A2(n2281), .B1(memory_REGFILE_WRITE_DATA[16]), 
        .B2(n3020), .ZN(n391) );
  buffd1 U1237 ( .I(n3005), .Z(n3025) );
  aoi22d1 U1238 ( .A1(n2932), .A2(n2282), .B1(n384), .B2(n3003), .ZN(n6877) );
  aoi22d1 U1239 ( .A1(n2870), .A2(n2838), .B1(n3027), .B2(
        memory_REGFILE_WRITE_DATA[17]), .ZN(n386) );
  aoi22d1 U1240 ( .A1(n3026), .A2(n388), .B1(n2984), .B2(
        memory_REGFILE_WRITE_DATA[15]), .ZN(n385) );
  oai211d1 U1241 ( .C1(n3025), .C2(n6877), .A(n386), .B(n385), .ZN(n387) );
  aon211d1 U1242 ( .C1(n3026), .C2(n2282), .B(n387), .A(n2856), .ZN(n390) );
  inv0d0 U1243 ( .I(CsrPlugin_mepc[15]), .ZN(n3611) );
  aoi22d1 U1244 ( .A1(n2328), .A2(_zz_CsrPlugin_csrMapping_readDataInit[15]), 
        .B1(n2327), .B2(CsrPlugin_mtval[15]), .ZN(n393) );
  oai21d1 U1245 ( .B1(n3611), .B2(n2541), .A(n393), .ZN(n2285) );
  aoi22d1 U1246 ( .A1(n2872), .A2(n2285), .B1(memory_REGFILE_WRITE_DATA[15]), 
        .B2(n3020), .ZN(n404) );
  inv0d0 U1247 ( .I(n2848), .ZN(n2284) );
  mx02d1 U1248 ( .I0(n2848), .I1(n2284), .S(n400), .Z(n3740) );
  aoi22d1 U1249 ( .A1(n2932), .A2(n2848), .B1(n396), .B2(n3003), .ZN(n6884) );
  aoi22d1 U1250 ( .A1(n2870), .A2(n2282), .B1(n3027), .B2(
        memory_REGFILE_WRITE_DATA[16]), .ZN(n398) );
  aoi22d1 U1251 ( .A1(n3026), .A2(n400), .B1(n2984), .B2(
        memory_REGFILE_WRITE_DATA[14]), .ZN(n397) );
  oai211d1 U1252 ( .C1(n3005), .C2(n6884), .A(n398), .B(n397), .ZN(n399) );
  aon211d1 U1253 ( .C1(n2960), .C2(n3740), .B(n399), .A(n2856), .ZN(n403) );
  aon211d1 U1254 ( .C1(n3040), .C2(n400), .B(n2989), .A(n2848), .ZN(n402) );
  nd02d0 U1255 ( .A1(n2923), .A2(n2863), .ZN(n401) );
  nd03d0 U1256 ( .A1(n405), .A2(_zz_lastStageRegFileWrite_payload_address_28), 
        .A3(_zz_lastStageRegFileWrite_payload_address_29), .ZN(n2393) );
  or02d2 U1257 ( .A1(\IBusCachedPlugin_cache/decodeStage_hit_valid ), .A2(
        n2359), .Z(n3049) );
  buffd1 U1258 ( .I(n3049), .Z(n3051) );
  nr02d0 U1259 ( .A1(n3050), .A2(n2214), .ZN(n2397) );
  inv0d0 U1260 ( .I(IBusCachedPlugin_fetchPc_booted), .ZN(n3287) );
  aoi211d1 U1261 ( .C1(n2374), .C2(n2397), .A(n3287), .B(reset), .ZN(n407) );
  inv0d0 U1262 ( .I(n407), .ZN(n2405) );
  nr02d1 U1263 ( .A1(n2393), .A2(n2405), .ZN(n454) );
  an03d1 U1264 ( .A1(n7121), .A2(IBusCachedPlugin_fetchPc_booted), .A3(n2399), 
        .Z(n525) );
  aoi22d1 U1265 ( .A1(n454), .A2(CsrPlugin_mepc[23]), .B1(n525), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[23]), .ZN(
        n410) );
  an02d1 U1266 ( .A1(n2397), .A2(n407), .Z(n544) );
  nr02d1 U1267 ( .A1(reset), .A2(n407), .ZN(n2382) );
  buffd1 U1268 ( .I(n2382), .Z(n540) );
  aoi22d1 U1269 ( .A1(n544), .A2(n406), .B1(n540), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[23]), .ZN(n409) );
  inv0d0 U1270 ( .I(n2393), .ZN(n2394) );
  nr02d0 U1271 ( .A1(n2137), .A2(n2367), .ZN(n2398) );
  an02d1 U1272 ( .A1(n2398), .A2(n407), .Z(n503) );
  aoi22d1 U1273 ( .A1(n531), .A2(CsrPlugin_mtvec_base[21]), .B1(n503), .B2(
        memory_BRANCH_CALC[23]), .ZN(n408) );
  aoi22d1 U1274 ( .A1(n454), .A2(CsrPlugin_mepc[26]), .B1(n525), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[26]), .ZN(
        n415) );
  buffd1 U1275 ( .I(n503), .Z(n542) );
  aoi22d1 U1276 ( .A1(n2382), .A2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[26]), .B1(n542), .B2(
        memory_BRANCH_CALC[26]), .ZN(n414) );
  buffd1 U1277 ( .I(n544), .Z(n534) );
  ah01d1 U1278 ( .A(n411), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[23]), .CO(n478), .S(
        n406) );
  aoi22d1 U1279 ( .A1(n531), .A2(CsrPlugin_mtvec_base[24]), .B1(n534), .B2(
        n412), .ZN(n413) );
  aoi22d1 U1280 ( .A1(n454), .A2(CsrPlugin_mepc[29]), .B1(n525), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[29]), .ZN(
        n421) );
  aoi22d1 U1281 ( .A1(n416), .A2(CsrPlugin_mtvec_base[27]), .B1(n542), .B2(
        memory_BRANCH_CALC[29]), .ZN(n420) );
  ah01d1 U1282 ( .A(n417), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[26]), .CO(n432), .S(
        n412) );
  aoi22d1 U1283 ( .A1(n534), .A2(n418), .B1(n2382), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[29]), .ZN(n419) );
  buffd1 U1284 ( .I(n525), .Z(n538) );
  aoi22d1 U1285 ( .A1(n538), .A2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[10]), .B1(
        n542), .B2(memory_BRANCH_CALC[10]), .ZN(n426) );
  aoi22d1 U1286 ( .A1(n416), .A2(CsrPlugin_mtvec_base[8]), .B1(n540), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[10]), .ZN(n425) );
  ah01d1 U1287 ( .A(n422), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[10]), .CO(n442), .S(
        n423) );
  aoi22d1 U1288 ( .A1(n454), .A2(CsrPlugin_mepc[10]), .B1(n534), .B2(n423), 
        .ZN(n424) );
  aoi22d1 U1289 ( .A1(n454), .A2(CsrPlugin_mepc[7]), .B1(n525), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[7]), .ZN(n431) );
  aoi22d1 U1290 ( .A1(n531), .A2(CsrPlugin_mtvec_base[5]), .B1(n542), .B2(
        memory_BRANCH_CALC[7]), .ZN(n430) );
  ah01d1 U1291 ( .A(n427), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[7]), .CO(n520), .S(
        n428) );
  aoi22d1 U1292 ( .A1(n534), .A2(n428), .B1(n2382), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[7]), .ZN(n429) );
  aoi22d1 U1293 ( .A1(n538), .A2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[27]), .B1(
        n540), .B2(IBusCachedPlugin_iBusRsp_stages_1_input_payload[27]), .ZN(
        n436) );
  aoi22d1 U1294 ( .A1(n531), .A2(CsrPlugin_mtvec_base[25]), .B1(n542), .B2(
        memory_BRANCH_CALC[27]), .ZN(n435) );
  ah01d1 U1295 ( .A(n432), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[27]), .CO(n532), .S(
        n433) );
  aoi22d1 U1296 ( .A1(n454), .A2(CsrPlugin_mepc[27]), .B1(n534), .B2(n433), 
        .ZN(n434) );
  aoi22d1 U1297 ( .A1(n531), .A2(CsrPlugin_mtvec_base[10]), .B1(n538), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[12]), .ZN(
        n441) );
  aoi22d1 U1298 ( .A1(n2382), .A2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[12]), .B1(n542), .B2(
        memory_BRANCH_CALC[12]), .ZN(n440) );
  ah01d1 U1299 ( .A(n437), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[12]), .CO(n447), .S(
        n438) );
  aoi22d1 U1300 ( .A1(n454), .A2(CsrPlugin_mepc[12]), .B1(n534), .B2(n438), 
        .ZN(n439) );
  aoi22d1 U1301 ( .A1(n531), .A2(CsrPlugin_mtvec_base[9]), .B1(n538), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[11]), .ZN(
        n446) );
  aoi22d1 U1302 ( .A1(n454), .A2(CsrPlugin_mepc[11]), .B1(n542), .B2(
        memory_BRANCH_CALC[11]), .ZN(n445) );
  ah01d1 U1303 ( .A(n442), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[11]), .CO(n437), .S(
        n443) );
  aoi22d1 U1304 ( .A1(n534), .A2(n443), .B1(n540), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[11]), .ZN(n444) );
  aoi22d1 U1305 ( .A1(n538), .A2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[13]), .B1(
        n540), .B2(IBusCachedPlugin_iBusRsp_stages_1_input_payload[13]), .ZN(
        n451) );
  ah01d1 U1306 ( .A(n447), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[13]), .CO(n541), .S(
        n448) );
  aoi22d1 U1307 ( .A1(n534), .A2(n448), .B1(n542), .B2(memory_BRANCH_CALC[13]), 
        .ZN(n450) );
  aoi22d1 U1308 ( .A1(n454), .A2(CsrPlugin_mepc[13]), .B1(n531), .B2(
        CsrPlugin_mtvec_base[11]), .ZN(n449) );
  ah01d1 U1309 ( .A(n452), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[6]), .CO(n427), .S(
        n453) );
  aoi22d1 U1310 ( .A1(n534), .A2(n453), .B1(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[6]), .B2(n538), .ZN(n457) );
  aoi22d1 U1311 ( .A1(IBusCachedPlugin_iBusRsp_stages_1_input_payload[6]), 
        .A2(n2382), .B1(memory_BRANCH_CALC[6]), .B2(n542), .ZN(n456) );
  buffd1 U1312 ( .I(n454), .Z(n539) );
  aoi22d1 U1313 ( .A1(CsrPlugin_mepc[6]), .A2(n539), .B1(
        CsrPlugin_mtvec_base[4]), .B2(n531), .ZN(n455) );
  aoi22d1 U1314 ( .A1(n538), .A2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[22]), .B1(
        n540), .B2(IBusCachedPlugin_iBusRsp_stages_1_input_payload[22]), .ZN(
        n462) );
  ah01d1 U1315 ( .A(n458), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[22]), .CO(n411), .S(
        n459) );
  aoi22d1 U1316 ( .A1(n544), .A2(n459), .B1(n503), .B2(memory_BRANCH_CALC[22]), 
        .ZN(n461) );
  aoi22d1 U1317 ( .A1(n539), .A2(CsrPlugin_mepc[22]), .B1(n531), .B2(
        CsrPlugin_mtvec_base[20]), .ZN(n460) );
  ah01d1 U1318 ( .A(n463), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[25]), .CO(n417), .S(
        n464) );
  aoi22d1 U1319 ( .A1(n544), .A2(n464), .B1(n538), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[25]), .ZN(
        n467) );
  aoi22d1 U1320 ( .A1(n416), .A2(CsrPlugin_mtvec_base[23]), .B1(n540), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[25]), .ZN(n466) );
  aoi22d1 U1321 ( .A1(n539), .A2(CsrPlugin_mepc[25]), .B1(n542), .B2(
        memory_BRANCH_CALC[25]), .ZN(n465) );
  ah01d1 U1322 ( .A(n468), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[18]), .CO(n510), .S(
        n469) );
  aoi22d1 U1323 ( .A1(n534), .A2(n469), .B1(n538), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[18]), .ZN(
        n472) );
  aoi22d1 U1324 ( .A1(n416), .A2(CsrPlugin_mtvec_base[16]), .B1(n540), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[18]), .ZN(n471) );
  aoi22d1 U1325 ( .A1(n539), .A2(CsrPlugin_mepc[18]), .B1(n503), .B2(
        memory_BRANCH_CALC[18]), .ZN(n470) );
  ah01d1 U1326 ( .A(n473), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[20]), .CO(n488), .S(
        n474) );
  aoi22d1 U1327 ( .A1(n544), .A2(n474), .B1(n525), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[20]), .ZN(
        n477) );
  aoi22d1 U1328 ( .A1(n539), .A2(CsrPlugin_mepc[20]), .B1(n503), .B2(
        memory_BRANCH_CALC[20]), .ZN(n476) );
  aoi22d1 U1329 ( .A1(n416), .A2(CsrPlugin_mtvec_base[18]), .B1(n540), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[20]), .ZN(n475) );
  aoi22d1 U1330 ( .A1(n531), .A2(CsrPlugin_mtvec_base[22]), .B1(n525), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[24]), .ZN(
        n482) );
  ah01d1 U1331 ( .A(n478), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[24]), .CO(n463), .S(
        n479) );
  aoi22d1 U1332 ( .A1(n544), .A2(n479), .B1(n503), .B2(memory_BRANCH_CALC[24]), 
        .ZN(n481) );
  aoi22d1 U1333 ( .A1(n539), .A2(CsrPlugin_mepc[24]), .B1(n540), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[24]), .ZN(n480) );
  ah01d1 U1334 ( .A(n483), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[17]), .CO(n468), .S(
        n484) );
  aoi22d1 U1335 ( .A1(n544), .A2(n484), .B1(n525), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[17]), .ZN(
        n487) );
  aoi22d1 U1336 ( .A1(n416), .A2(CsrPlugin_mtvec_base[15]), .B1(n503), .B2(
        memory_BRANCH_CALC[17]), .ZN(n486) );
  aoi22d1 U1337 ( .A1(n539), .A2(CsrPlugin_mepc[17]), .B1(n540), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[17]), .ZN(n485) );
  aoi22d1 U1338 ( .A1(n538), .A2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[21]), .B1(
        n503), .B2(memory_BRANCH_CALC[21]), .ZN(n492) );
  ah01d1 U1339 ( .A(n488), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[21]), .CO(n458), .S(
        n489) );
  aoi22d1 U1340 ( .A1(n416), .A2(CsrPlugin_mtvec_base[19]), .B1(n534), .B2(
        n489), .ZN(n491) );
  aoi22d1 U1341 ( .A1(n539), .A2(CsrPlugin_mepc[21]), .B1(n540), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[21]), .ZN(n490) );
  aoi22d1 U1342 ( .A1(n538), .A2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[15]), .B1(
        n503), .B2(memory_BRANCH_CALC[15]), .ZN(n497) );
  aoi22d1 U1343 ( .A1(n531), .A2(CsrPlugin_mtvec_base[13]), .B1(n540), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[15]), .ZN(n496) );
  ah01d1 U1344 ( .A(n493), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[15]), .CO(n526), .S(
        n494) );
  aoi22d1 U1345 ( .A1(n539), .A2(CsrPlugin_mepc[15]), .B1(n534), .B2(n494), 
        .ZN(n495) );
  aoi22d1 U1346 ( .A1(n531), .A2(CsrPlugin_mtvec_base[7]), .B1(n538), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[9]), .ZN(n502) );
  aoi22d1 U1347 ( .A1(n2382), .A2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[9]), .B1(n542), .B2(
        memory_BRANCH_CALC[9]), .ZN(n501) );
  ah01d1 U1348 ( .A(n498), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[9]), .CO(n422), .S(
        n499) );
  aoi22d1 U1349 ( .A1(n539), .A2(CsrPlugin_mepc[9]), .B1(n534), .B2(n499), 
        .ZN(n500) );
  aoi22d1 U1350 ( .A1(n531), .A2(CsrPlugin_mtvec_base[29]), .B1(n525), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[31]), .ZN(
        n509) );
  aoi22d1 U1351 ( .A1(n539), .A2(CsrPlugin_mepc[31]), .B1(n503), .B2(
        memory_BRANCH_CALC[31]), .ZN(n508) );
  ah01d1 U1352 ( .A(n504), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[29]), .CO(n515), .S(
        n418) );
  xr02d1 U1353 ( .A1(n505), .A2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[31]), .Z(n506) );
  aoi22d1 U1354 ( .A1(n544), .A2(n506), .B1(n540), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[31]), .ZN(n507) );
  aoi22d1 U1355 ( .A1(n538), .A2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[19]), .B1(
        n540), .B2(IBusCachedPlugin_iBusRsp_stages_1_input_payload[19]), .ZN(
        n514) );
  aoi22d1 U1356 ( .A1(n539), .A2(CsrPlugin_mepc[19]), .B1(n531), .B2(
        CsrPlugin_mtvec_base[17]), .ZN(n513) );
  ah01d1 U1357 ( .A(n510), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[19]), .CO(n473), .S(
        n511) );
  aoi22d1 U1358 ( .A1(n534), .A2(n511), .B1(n542), .B2(memory_BRANCH_CALC[19]), 
        .ZN(n512) );
  aoi22d1 U1359 ( .A1(n416), .A2(CsrPlugin_mtvec_base[28]), .B1(n538), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[30]), .ZN(
        n519) );
  ah01d1 U1360 ( .A(n515), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[30]), .CO(n505), .S(
        n516) );
  aoi22d1 U1361 ( .A1(n544), .A2(n516), .B1(n542), .B2(memory_BRANCH_CALC[30]), 
        .ZN(n518) );
  aoi22d1 U1362 ( .A1(n539), .A2(CsrPlugin_mepc[30]), .B1(n2382), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[30]), .ZN(n517) );
  aoi22d1 U1363 ( .A1(n531), .A2(CsrPlugin_mtvec_base[6]), .B1(n538), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[8]), .ZN(n524) );
  ah01d1 U1364 ( .A(n520), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[8]), .CO(n498), .S(
        n521) );
  aoi22d1 U1365 ( .A1(n539), .A2(CsrPlugin_mepc[8]), .B1(n534), .B2(n521), 
        .ZN(n523) );
  aoi22d1 U1366 ( .A1(n2382), .A2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[8]), .B1(n542), .B2(
        memory_BRANCH_CALC[8]), .ZN(n522) );
  aoi22d1 U1367 ( .A1(n539), .A2(CsrPlugin_mepc[16]), .B1(n525), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[16]), .ZN(
        n530) );
  ah01d1 U1368 ( .A(n526), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[16]), .CO(n483), .S(
        n527) );
  aoi22d1 U1369 ( .A1(n534), .A2(n527), .B1(n542), .B2(memory_BRANCH_CALC[16]), 
        .ZN(n529) );
  aoi22d1 U1370 ( .A1(n531), .A2(CsrPlugin_mtvec_base[14]), .B1(n540), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[16]), .ZN(n528) );
  aoi22d1 U1371 ( .A1(n531), .A2(CsrPlugin_mtvec_base[26]), .B1(n538), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[28]), .ZN(
        n537) );
  aoi22d1 U1372 ( .A1(n539), .A2(CsrPlugin_mepc[28]), .B1(n2382), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[28]), .ZN(n536) );
  ah01d1 U1373 ( .A(n532), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[28]), .CO(n504), .S(
        n533) );
  aoi22d1 U1374 ( .A1(n534), .A2(n533), .B1(n542), .B2(memory_BRANCH_CALC[28]), 
        .ZN(n535) );
  aoi22d1 U1375 ( .A1(n539), .A2(CsrPlugin_mepc[14]), .B1(n538), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[14]), .ZN(
        n547) );
  aoi22d1 U1376 ( .A1(n531), .A2(CsrPlugin_mtvec_base[12]), .B1(n540), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[14]), .ZN(n546) );
  ah01d1 U1377 ( .A(n541), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[14]), .CO(n493), .S(
        n543) );
  aoi22d1 U1378 ( .A1(n544), .A2(n543), .B1(n542), .B2(memory_BRANCH_CALC[14]), 
        .ZN(n545) );
  nr02d0 U1379 ( .A1(n6977), .A2(n556), .ZN(n555) );
  aoi22d1 U1380 ( .A1(dBusWishbone_CYC), .A2(dBusWishbone_DAT_MOSI[10]), .B1(
        execute_RS2[10]), .B2(n555), .ZN(n548) );
  inv0d2 U1381 ( .I(n6977), .ZN(n6963) );
  nd03d0 U1382 ( .A1(n556), .A2(execute_RS2[2]), .A3(n6963), .ZN(n6978) );
  nd02d0 U1383 ( .A1(n548), .A2(n6978), .ZN(n3872) );
  aoi22d1 U1384 ( .A1(dBusWishbone_CYC), .A2(dBusWishbone_DAT_MOSI[9]), .B1(
        execute_RS2[9]), .B2(n555), .ZN(n549) );
  inv0d0 U1385 ( .I(dBusWishbone_CYC), .ZN(n6920) );
  nd03d0 U1386 ( .A1(n556), .A2(execute_RS2[1]), .A3(n6920), .ZN(n6989) );
  nd02d0 U1387 ( .A1(n549), .A2(n6989), .ZN(n3867) );
  aoi22d1 U1388 ( .A1(dBusWishbone_CYC), .A2(dBusWishbone_DAT_MOSI[13]), .B1(
        execute_RS2[13]), .B2(n555), .ZN(n550) );
  nd03d0 U1389 ( .A1(n556), .A2(execute_RS2[5]), .A3(n6963), .ZN(n6953) );
  nd02d0 U1390 ( .A1(n550), .A2(n6953), .ZN(n3887) );
  aoi22d1 U1391 ( .A1(n6977), .A2(dBusWishbone_DAT_MOSI[14]), .B1(
        execute_RS2[14]), .B2(n555), .ZN(n551) );
  nd03d0 U1392 ( .A1(n556), .A2(execute_RS2[6]), .A3(n6963), .ZN(n6946) );
  nd02d0 U1393 ( .A1(n551), .A2(n6946), .ZN(n3892) );
  aoi22d1 U1394 ( .A1(n6977), .A2(dBusWishbone_DAT_MOSI[8]), .B1(
        execute_RS2[8]), .B2(n555), .ZN(n552) );
  nd03d0 U1395 ( .A1(n556), .A2(execute_RS2[0]), .A3(n6963), .ZN(n6921) );
  nd02d0 U1396 ( .A1(n552), .A2(n6921), .ZN(n3905) );
  aoi22d1 U1397 ( .A1(n6977), .A2(dBusWishbone_DAT_MOSI[15]), .B1(
        execute_RS2[15]), .B2(n555), .ZN(n553) );
  nd03d0 U1398 ( .A1(n556), .A2(execute_RS2[7]), .A3(n6963), .ZN(n6933) );
  nd02d0 U1399 ( .A1(n553), .A2(n6933), .ZN(n3899) );
  aoi22d1 U1400 ( .A1(dBusWishbone_CYC), .A2(dBusWishbone_DAT_MOSI[11]), .B1(
        execute_RS2[11]), .B2(n555), .ZN(n554) );
  nd03d0 U1401 ( .A1(n556), .A2(execute_RS2[3]), .A3(n6963), .ZN(n6969) );
  nd02d0 U1402 ( .A1(n554), .A2(n6969), .ZN(n3877) );
  aoi22d1 U1403 ( .A1(dBusWishbone_CYC), .A2(dBusWishbone_DAT_MOSI[12]), .B1(
        execute_RS2[12]), .B2(n555), .ZN(n557) );
  inv0d1 U1404 ( .I(n6977), .ZN(n6972) );
  nd03d0 U1405 ( .A1(n556), .A2(execute_RS2[4]), .A3(n6972), .ZN(n6960) );
  nd02d0 U1406 ( .A1(n557), .A2(n6960), .ZN(n3882) );
  inv0d1 U1407 ( .I(n2193), .ZN(n2209) );
  aoi22d1 U1408 ( .A1(execute_INSTRUCTION[0]), .A2(n2209), .B1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[0]), .B2(n2181), 
        .ZN(n560) );
  buffd1 U1409 ( .I(n2190), .Z(n2186) );
  aoi22d1 U1410 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[0]), .A2(n2186), .B1(
        n2198), .B2(memory_REGFILE_WRITE_DATA[0]), .ZN(n559) );
  nd02d0 U1411 ( .A1(n560), .A2(n559), .ZN(n6207) );
  an02d0 U1412 ( .A1(n561), .A2(CsrPlugin_pipelineLiberator_pcValids_1), .Z(
        n6133) );
  inv0d0 U1413 ( .I(execute_CSR_WRITE_OPCODE), .ZN(n2551) );
  aoi21d1 U1414 ( .B1(_zz__zz_execute_BranchPlugin_branch_src2[12]), .B2(n564), 
        .A(n563), .ZN(n565) );
  aoim21d1 U1415 ( .B1(n2289), .B2(n3008), .A(n565), .ZN(n2349) );
  an03d0 U1416 ( .A1(n3566), .A2(execute_CsrPlugin_csr_836), .A3(n2349), .Z(
        N2007) );
  inv0d0 U1417 ( .I(IBusCachedPlugin_cache_io_cpu_fetch_data[15]), .ZN(n6636)
         );
  mx02d1 U1418 ( .I0(n6636), .I1(n174), .S(n2374), .Z(n571) );
  mx02d1 U1419 ( .I0(IBusCachedPlugin_cache_io_cpu_fetch_data[16]), .I1(
        decode_INSTRUCTION[16]), .S(n2374), .Z(n569) );
  inv0d0 U1420 ( .I(IBusCachedPlugin_cache_io_cpu_fetch_data[17]), .ZN(n6611)
         );
  mx02d1 U1421 ( .I0(n6611), .I1(n2622), .S(n2374), .Z(n580) );
  inv0d0 U1422 ( .I(IBusCachedPlugin_cache_io_cpu_fetch_data[19]), .ZN(n6586)
         );
  mx02d1 U1423 ( .I0(n6586), .I1(n2618), .S(n2374), .Z(n567) );
  inv0d0 U1424 ( .I(IBusCachedPlugin_cache_io_cpu_fetch_data[18]), .ZN(n6598)
         );
  mx02d1 U1425 ( .I0(n6598), .I1(n173), .S(n2374), .Z(n566) );
  nr02d0 U1426 ( .A1(n567), .A2(n566), .ZN(n583) );
  nr02d1 U1427 ( .A1(n590), .A2(n589), .ZN(n1138) );
  buffd1 U1428 ( .I(n1138), .Z(n1195) );
  inv0d0 U1429 ( .I(n569), .ZN(n572) );
  inv0d0 U1430 ( .I(n571), .ZN(n568) );
  inv0d0 U1431 ( .I(n567), .ZN(n579) );
  nr02d0 U1432 ( .A1(n566), .A2(n579), .ZN(n573) );
  inv0d0 U1433 ( .I(n580), .ZN(n582) );
  nr02d1 U1434 ( .A1(n597), .A2(n595), .ZN(n1072) );
  buffd1 U1435 ( .I(n1072), .Z(n1244) );
  aoi22d1 U1436 ( .A1(\RegFilePlugin_regFile[26][31] ), .A2(n1195), .B1(
        \RegFilePlugin_regFile[13][31] ), .B2(n1244), .ZN(n577) );
  inv0d0 U1437 ( .I(n566), .ZN(n578) );
  nr02d0 U1438 ( .A1(n567), .A2(n578), .ZN(n570) );
  nr02d1 U1439 ( .A1(n597), .A2(n601), .ZN(n1099) );
  buffd1 U1440 ( .I(n1099), .Z(n1251) );
  buffd1 U1441 ( .I(n758), .Z(n1190) );
  aoi22d1 U1442 ( .A1(\RegFilePlugin_regFile[17][31] ), .A2(n1251), .B1(
        \RegFilePlugin_regFile[19][31] ), .B2(n1190), .ZN(n576) );
  nr02d1 U1443 ( .A1(n599), .A2(n600), .ZN(n889) );
  buffd1 U1444 ( .I(n889), .Z(n1222) );
  buffd1 U1445 ( .I(n1185), .Z(n1294) );
  aoi22d1 U1446 ( .A1(\RegFilePlugin_regFile[20][31] ), .A2(n1222), .B1(
        \RegFilePlugin_regFile[8][31] ), .B2(n1294), .ZN(n575) );
  nr02d1 U1447 ( .A1(n589), .A2(n597), .ZN(n842) );
  buffd1 U1448 ( .I(n842), .Z(n1148) );
  buffd1 U1449 ( .I(n736), .Z(n1282) );
  aoi22d1 U1450 ( .A1(\RegFilePlugin_regFile[25][31] ), .A2(n1148), .B1(
        \RegFilePlugin_regFile[14][31] ), .B2(n1282), .ZN(n574) );
  nr02d0 U1451 ( .A1(n579), .A2(n578), .ZN(n581) );
  nr02d1 U1452 ( .A1(n590), .A2(n596), .ZN(n1073) );
  nr02d1 U1453 ( .A1(n590), .A2(n599), .ZN(n1143) );
  buffd1 U1454 ( .I(n1143), .Z(n1288) );
  aoi22d1 U1455 ( .A1(\RegFilePlugin_regFile[2][31] ), .A2(n1073), .B1(
        \RegFilePlugin_regFile[22][31] ), .B2(n1288), .ZN(n587) );
  buffd1 U1456 ( .I(n699), .Z(n1269) );
  nr02d1 U1457 ( .A1(n590), .A2(n598), .ZN(n658) );
  buffd1 U1458 ( .I(n658), .Z(n1208) );
  aoi22d1 U1459 ( .A1(\RegFilePlugin_regFile[1][31] ), .A2(n1269), .B1(
        \RegFilePlugin_regFile[10][31] ), .B2(n1208), .ZN(n586) );
  buffd1 U1460 ( .I(n1216), .Z(n1253) );
  nr02d1 U1461 ( .A1(n590), .A2(n602), .ZN(n653) );
  buffd1 U1462 ( .I(n653), .Z(n1260) );
  aoi22d1 U1463 ( .A1(\RegFilePlugin_regFile[7][31] ), .A2(n1253), .B1(
        \RegFilePlugin_regFile[30][31] ), .B2(n1260), .ZN(n585) );
  nr02d1 U1464 ( .A1(n597), .A2(n588), .ZN(n757) );
  buffd1 U1465 ( .I(n757), .Z(n1166) );
  nr02d1 U1466 ( .A1(n600), .A2(n588), .ZN(n1238) );
  buffd1 U1467 ( .I(n1238), .Z(n1217) );
  aoi22d1 U1468 ( .A1(\RegFilePlugin_regFile[5][31] ), .A2(n1166), .B1(
        \RegFilePlugin_regFile[4][31] ), .B2(n1217), .ZN(n584) );
  nr02d1 U1469 ( .A1(n597), .A2(n602), .ZN(n1094) );
  buffd1 U1470 ( .I(n1094), .Z(n1271) );
  nr02d1 U1471 ( .A1(n603), .A2(n596), .ZN(n1210) );
  buffd1 U1472 ( .I(n1210), .Z(n1280) );
  aoi22d1 U1473 ( .A1(\RegFilePlugin_regFile[29][31] ), .A2(n1271), .B1(
        \RegFilePlugin_regFile[3][31] ), .B2(n1280), .ZN(n594) );
  buffd1 U1474 ( .I(n1161), .Z(n1250) );
  nr02d1 U1475 ( .A1(n595), .A2(n603), .ZN(n1116) );
  buffd1 U1476 ( .I(n1116), .Z(n1209) );
  aoi22d1 U1477 ( .A1(\RegFilePlugin_regFile[6][31] ), .A2(n1250), .B1(
        \RegFilePlugin_regFile[15][31] ), .B2(n1209), .ZN(n593) );
  nr02d1 U1478 ( .A1(n600), .A2(n602), .ZN(n988) );
  buffd1 U1479 ( .I(n988), .Z(n1298) );
  nr02d1 U1480 ( .A1(n589), .A2(n600), .ZN(n867) );
  aoi22d1 U1481 ( .A1(\RegFilePlugin_regFile[28][31] ), .A2(n1298), .B1(
        \RegFilePlugin_regFile[24][31] ), .B2(n867), .ZN(n592) );
  buffd1 U1482 ( .I(n780), .Z(n1270) );
  buffd1 U1483 ( .I(n612), .Z(n1297) );
  aoi22d1 U1484 ( .A1(\RegFilePlugin_regFile[27][31] ), .A2(n1270), .B1(
        \RegFilePlugin_regFile[18][31] ), .B2(n1297), .ZN(n591) );
  nr02d1 U1485 ( .A1(n595), .A2(n600), .ZN(n884) );
  buffd1 U1486 ( .I(n884), .Z(n1296) );
  buffd1 U1487 ( .I(n987), .Z(n1258) );
  aoi22d1 U1488 ( .A1(\RegFilePlugin_regFile[12][31] ), .A2(n1296), .B1(
        \RegFilePlugin_regFile[21][31] ), .B2(n1258), .ZN(n607) );
  nr02d1 U1489 ( .A1(n600), .A2(n596), .ZN(n926) );
  buffd1 U1490 ( .I(n926), .Z(n1215) );
  nr02d1 U1491 ( .A1(n597), .A2(n598), .ZN(n841) );
  buffd1 U1492 ( .I(n841), .Z(n1229) );
  aoi22d1 U1493 ( .A1(\RegFilePlugin_regFile[0][31] ), .A2(n1215), .B1(
        \RegFilePlugin_regFile[9][31] ), .B2(n1229), .ZN(n606) );
  buffd1 U1494 ( .I(n989), .Z(n1171) );
  nr02d1 U1495 ( .A1(n603), .A2(n599), .ZN(n779) );
  buffd1 U1496 ( .I(n779), .Z(n1281) );
  aoi22d1 U1497 ( .A1(\RegFilePlugin_regFile[11][31] ), .A2(n1171), .B1(
        \RegFilePlugin_regFile[23][31] ), .B2(n1281), .ZN(n605) );
  nr02d1 U1498 ( .A1(n601), .A2(n600), .ZN(n1010) );
  buffd1 U1499 ( .I(n1010), .Z(n1274) );
  nr02d1 U1500 ( .A1(n603), .A2(n602), .ZN(n1011) );
  buffd1 U1501 ( .I(n1011), .Z(n1228) );
  aoi22d1 U1502 ( .A1(\RegFilePlugin_regFile[16][31] ), .A2(n1274), .B1(
        \RegFilePlugin_regFile[31][31] ), .B2(n1228), .ZN(n604) );
  or04d0 U1503 ( .A1(n611), .A2(n610), .A3(n609), .A4(n608), .Z(N823) );
  buffd1 U1504 ( .I(n612), .Z(n1223) );
  aoi22d1 U1505 ( .A1(n1210), .A2(\RegFilePlugin_regFile[3][28] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][28] ), .ZN(n616) );
  aoi22d1 U1506 ( .A1(n926), .A2(\RegFilePlugin_regFile[0][28] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][28] ), .ZN(n615) );
  aoi22d1 U1507 ( .A1(n889), .A2(\RegFilePlugin_regFile[20][28] ), .B1(n884), 
        .B2(\RegFilePlugin_regFile[12][28] ), .ZN(n614) );
  aoi22d1 U1508 ( .A1(n1073), .A2(\RegFilePlugin_regFile[2][28] ), .B1(n1208), 
        .B2(\RegFilePlugin_regFile[10][28] ), .ZN(n613) );
  aoi22d1 U1509 ( .A1(n1260), .A2(\RegFilePlugin_regFile[30][28] ), .B1(n757), 
        .B2(\RegFilePlugin_regFile[5][28] ), .ZN(n620) );
  aoi22d1 U1510 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][28] ), .B1(n988), 
        .B2(\RegFilePlugin_regFile[28][28] ), .ZN(n619) );
  buffd1 U1511 ( .I(n1185), .Z(n1239) );
  aoi22d1 U1512 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][28] ), .B1(n842), 
        .B2(\RegFilePlugin_regFile[25][28] ), .ZN(n618) );
  aoi22d1 U1513 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][28] ), .B1(n1190), 
        .B2(\RegFilePlugin_regFile[19][28] ), .ZN(n617) );
  buffd1 U1514 ( .I(n989), .Z(n1272) );
  aoi22d1 U1515 ( .A1(n1272), .A2(\RegFilePlugin_regFile[11][28] ), .B1(n1281), 
        .B2(\RegFilePlugin_regFile[23][28] ), .ZN(n624) );
  aoi22d1 U1516 ( .A1(n1271), .A2(\RegFilePlugin_regFile[29][28] ), .B1(n867), 
        .B2(\RegFilePlugin_regFile[24][28] ), .ZN(n623) );
  buffd1 U1517 ( .I(n987), .Z(n1295) );
  aoi22d1 U1518 ( .A1(n1295), .A2(\RegFilePlugin_regFile[21][28] ), .B1(n841), 
        .B2(\RegFilePlugin_regFile[9][28] ), .ZN(n622) );
  aoi22d1 U1519 ( .A1(n1072), .A2(\RegFilePlugin_regFile[13][28] ), .B1(n1282), 
        .B2(\RegFilePlugin_regFile[14][28] ), .ZN(n621) );
  buffd1 U1520 ( .I(n1216), .Z(n1289) );
  buffd1 U1521 ( .I(n1161), .Z(n1275) );
  aoi22d1 U1522 ( .A1(n1289), .A2(\RegFilePlugin_regFile[7][28] ), .B1(n1275), 
        .B2(\RegFilePlugin_regFile[6][28] ), .ZN(n628) );
  aoi22d1 U1523 ( .A1(n1269), .A2(\RegFilePlugin_regFile[1][28] ), .B1(n1270), 
        .B2(\RegFilePlugin_regFile[27][28] ), .ZN(n627) );
  aoi22d1 U1524 ( .A1(n1288), .A2(\RegFilePlugin_regFile[22][28] ), .B1(n1010), 
        .B2(\RegFilePlugin_regFile[16][28] ), .ZN(n626) );
  aoi22d1 U1525 ( .A1(n1217), .A2(\RegFilePlugin_regFile[4][28] ), .B1(n1209), 
        .B2(\RegFilePlugin_regFile[15][28] ), .ZN(n625) );
  or04d0 U1526 ( .A1(n632), .A2(n631), .A3(n630), .A4(n629), .Z(N826) );
  buffd1 U1527 ( .I(n699), .Z(n1259) );
  aoi22d1 U1528 ( .A1(n1259), .A2(\RegFilePlugin_regFile[1][26] ), .B1(n1209), 
        .B2(\RegFilePlugin_regFile[15][26] ), .ZN(n636) );
  aoi22d1 U1529 ( .A1(n658), .A2(\RegFilePlugin_regFile[10][26] ), .B1(n841), 
        .B2(\RegFilePlugin_regFile[9][26] ), .ZN(n635) );
  aoi22d1 U1530 ( .A1(n1288), .A2(\RegFilePlugin_regFile[22][26] ), .B1(n1210), 
        .B2(\RegFilePlugin_regFile[3][26] ), .ZN(n634) );
  aoi22d1 U1531 ( .A1(n1099), .A2(\RegFilePlugin_regFile[17][26] ), .B1(n757), 
        .B2(\RegFilePlugin_regFile[5][26] ), .ZN(n633) );
  aoi22d1 U1532 ( .A1(n1217), .A2(\RegFilePlugin_regFile[4][26] ), .B1(n1094), 
        .B2(\RegFilePlugin_regFile[29][26] ), .ZN(n640) );
  aoi22d1 U1533 ( .A1(n842), .A2(\RegFilePlugin_regFile[25][26] ), .B1(n653), 
        .B2(\RegFilePlugin_regFile[30][26] ), .ZN(n639) );
  aoi22d1 U1534 ( .A1(n1138), .A2(\RegFilePlugin_regFile[26][26] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][26] ), .ZN(n638) );
  aoi22d1 U1535 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][26] ), .B1(n1275), 
        .B2(\RegFilePlugin_regFile[6][26] ), .ZN(n637) );
  aoi22d1 U1536 ( .A1(n1072), .A2(\RegFilePlugin_regFile[13][26] ), .B1(n1171), 
        .B2(\RegFilePlugin_regFile[11][26] ), .ZN(n644) );
  buffd1 U1537 ( .I(n758), .Z(n1287) );
  aoi22d1 U1538 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][26] ), .B1(n1281), 
        .B2(\RegFilePlugin_regFile[23][26] ), .ZN(n643) );
  buffd1 U1539 ( .I(n1073), .Z(n1176) );
  aoi22d1 U1540 ( .A1(n1176), .A2(\RegFilePlugin_regFile[2][26] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][26] ), .ZN(n642) );
  buffd1 U1541 ( .I(n867), .Z(n1273) );
  aoi22d1 U1542 ( .A1(n1222), .A2(\RegFilePlugin_regFile[20][26] ), .B1(n1273), 
        .B2(\RegFilePlugin_regFile[24][26] ), .ZN(n641) );
  aoi22d1 U1543 ( .A1(n1289), .A2(\RegFilePlugin_regFile[7][26] ), .B1(n1010), 
        .B2(\RegFilePlugin_regFile[16][26] ), .ZN(n648) );
  aoi22d1 U1544 ( .A1(n1282), .A2(\RegFilePlugin_regFile[14][26] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][26] ), .ZN(n647) );
  aoi22d1 U1545 ( .A1(n1270), .A2(\RegFilePlugin_regFile[27][26] ), .B1(n1296), 
        .B2(\RegFilePlugin_regFile[12][26] ), .ZN(n646) );
  aoi22d1 U1546 ( .A1(n1298), .A2(\RegFilePlugin_regFile[28][26] ), .B1(n1258), 
        .B2(\RegFilePlugin_regFile[21][26] ), .ZN(n645) );
  or04d0 U1547 ( .A1(n652), .A2(n651), .A3(n650), .A4(n649), .Z(N828) );
  aoi22d1 U1548 ( .A1(n1244), .A2(\RegFilePlugin_regFile[13][27] ), .B1(n1259), 
        .B2(\RegFilePlugin_regFile[1][27] ), .ZN(n657) );
  aoi22d1 U1549 ( .A1(n1217), .A2(\RegFilePlugin_regFile[4][27] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][27] ), .ZN(n656) );
  aoi22d1 U1550 ( .A1(n1280), .A2(\RegFilePlugin_regFile[3][27] ), .B1(n1298), 
        .B2(\RegFilePlugin_regFile[28][27] ), .ZN(n655) );
  aoi22d1 U1551 ( .A1(n653), .A2(\RegFilePlugin_regFile[30][27] ), .B1(n1166), 
        .B2(\RegFilePlugin_regFile[5][27] ), .ZN(n654) );
  aoi22d1 U1552 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][27] ), .B1(n1171), 
        .B2(\RegFilePlugin_regFile[11][27] ), .ZN(n662) );
  aoi22d1 U1553 ( .A1(n1148), .A2(\RegFilePlugin_regFile[25][27] ), .B1(n658), 
        .B2(\RegFilePlugin_regFile[10][27] ), .ZN(n661) );
  aoi22d1 U1554 ( .A1(n1296), .A2(\RegFilePlugin_regFile[12][27] ), .B1(n1281), 
        .B2(\RegFilePlugin_regFile[23][27] ), .ZN(n660) );
  aoi22d1 U1555 ( .A1(n1176), .A2(\RegFilePlugin_regFile[2][27] ), .B1(n1010), 
        .B2(\RegFilePlugin_regFile[16][27] ), .ZN(n659) );
  aoi22d1 U1556 ( .A1(n1222), .A2(\RegFilePlugin_regFile[20][27] ), .B1(n1209), 
        .B2(\RegFilePlugin_regFile[15][27] ), .ZN(n666) );
  aoi22d1 U1557 ( .A1(n1271), .A2(\RegFilePlugin_regFile[29][27] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][27] ), .ZN(n665) );
  aoi22d1 U1558 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][27] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][27] ), .ZN(n664) );
  aoi22d1 U1559 ( .A1(n1275), .A2(\RegFilePlugin_regFile[6][27] ), .B1(n867), 
        .B2(\RegFilePlugin_regFile[24][27] ), .ZN(n663) );
  aoi22d1 U1560 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][27] ), .B1(n1258), 
        .B2(\RegFilePlugin_regFile[21][27] ), .ZN(n670) );
  aoi22d1 U1561 ( .A1(n1282), .A2(\RegFilePlugin_regFile[14][27] ), .B1(n1288), 
        .B2(\RegFilePlugin_regFile[22][27] ), .ZN(n669) );
  aoi22d1 U1562 ( .A1(n1289), .A2(\RegFilePlugin_regFile[7][27] ), .B1(n841), 
        .B2(\RegFilePlugin_regFile[9][27] ), .ZN(n668) );
  buffd1 U1563 ( .I(n780), .Z(n1252) );
  aoi22d1 U1564 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][27] ), .B1(n1252), 
        .B2(\RegFilePlugin_regFile[27][27] ), .ZN(n667) );
  or04d0 U1565 ( .A1(n674), .A2(n673), .A3(n672), .A4(n671), .Z(N827) );
  aoi22d1 U1566 ( .A1(n1217), .A2(\RegFilePlugin_regFile[4][25] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][25] ), .ZN(n678) );
  aoi22d1 U1567 ( .A1(n1260), .A2(\RegFilePlugin_regFile[30][25] ), .B1(n1010), 
        .B2(\RegFilePlugin_regFile[16][25] ), .ZN(n677) );
  aoi22d1 U1568 ( .A1(n1148), .A2(\RegFilePlugin_regFile[25][25] ), .B1(n1094), 
        .B2(\RegFilePlugin_regFile[29][25] ), .ZN(n676) );
  aoi22d1 U1569 ( .A1(n1222), .A2(\RegFilePlugin_regFile[20][25] ), .B1(n1281), 
        .B2(\RegFilePlugin_regFile[23][25] ), .ZN(n675) );
  aoi22d1 U1570 ( .A1(n1099), .A2(\RegFilePlugin_regFile[17][25] ), .B1(n841), 
        .B2(\RegFilePlugin_regFile[9][25] ), .ZN(n682) );
  aoi22d1 U1571 ( .A1(n1138), .A2(\RegFilePlugin_regFile[26][25] ), .B1(n1244), 
        .B2(\RegFilePlugin_regFile[13][25] ), .ZN(n681) );
  aoi22d1 U1572 ( .A1(n1208), .A2(\RegFilePlugin_regFile[10][25] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][25] ), .ZN(n680) );
  aoi22d1 U1573 ( .A1(n1166), .A2(\RegFilePlugin_regFile[5][25] ), .B1(n1275), 
        .B2(\RegFilePlugin_regFile[6][25] ), .ZN(n679) );
  aoi22d1 U1574 ( .A1(n988), .A2(\RegFilePlugin_regFile[28][25] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][25] ), .ZN(n686) );
  aoi22d1 U1575 ( .A1(n1176), .A2(\RegFilePlugin_regFile[2][25] ), .B1(n1273), 
        .B2(\RegFilePlugin_regFile[24][25] ), .ZN(n685) );
  aoi22d1 U1576 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][25] ), .B1(n1253), 
        .B2(\RegFilePlugin_regFile[7][25] ), .ZN(n684) );
  aoi22d1 U1577 ( .A1(n1282), .A2(\RegFilePlugin_regFile[14][25] ), .B1(n1209), 
        .B2(\RegFilePlugin_regFile[15][25] ), .ZN(n683) );
  aoi22d1 U1578 ( .A1(n1288), .A2(\RegFilePlugin_regFile[22][25] ), .B1(n1280), 
        .B2(\RegFilePlugin_regFile[3][25] ), .ZN(n690) );
  aoi22d1 U1579 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][25] ), .B1(n1296), 
        .B2(\RegFilePlugin_regFile[12][25] ), .ZN(n689) );
  aoi22d1 U1580 ( .A1(n1252), .A2(\RegFilePlugin_regFile[27][25] ), .B1(n1171), 
        .B2(\RegFilePlugin_regFile[11][25] ), .ZN(n688) );
  aoi22d1 U1581 ( .A1(n1259), .A2(\RegFilePlugin_regFile[1][25] ), .B1(n1258), 
        .B2(\RegFilePlugin_regFile[21][25] ), .ZN(n687) );
  or04d0 U1582 ( .A1(n694), .A2(n693), .A3(n692), .A4(n691), .Z(N829) );
  aoi22d1 U1583 ( .A1(n1238), .A2(\RegFilePlugin_regFile[4][11] ), .B1(n1010), 
        .B2(\RegFilePlugin_regFile[16][11] ), .ZN(n698) );
  buffd1 U1584 ( .I(n736), .Z(n1245) );
  aoi22d1 U1585 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][11] ), .B1(n1296), 
        .B2(\RegFilePlugin_regFile[12][11] ), .ZN(n697) );
  aoi22d1 U1586 ( .A1(n653), .A2(\RegFilePlugin_regFile[30][11] ), .B1(n1298), 
        .B2(\RegFilePlugin_regFile[28][11] ), .ZN(n696) );
  aoi22d1 U1587 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][11] ), .B1(n1288), 
        .B2(\RegFilePlugin_regFile[22][11] ), .ZN(n695) );
  aoi22d1 U1588 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][11] ), .B1(n1210), 
        .B2(\RegFilePlugin_regFile[3][11] ), .ZN(n703) );
  aoi22d1 U1589 ( .A1(n1244), .A2(\RegFilePlugin_regFile[13][11] ), .B1(n1270), 
        .B2(\RegFilePlugin_regFile[27][11] ), .ZN(n702) );
  aoi22d1 U1590 ( .A1(n699), .A2(\RegFilePlugin_regFile[1][11] ), .B1(n1273), 
        .B2(\RegFilePlugin_regFile[24][11] ), .ZN(n701) );
  aoi22d1 U1591 ( .A1(n1295), .A2(\RegFilePlugin_regFile[21][11] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][11] ), .ZN(n700) );
  aoi22d1 U1592 ( .A1(n1190), .A2(\RegFilePlugin_regFile[19][11] ), .B1(n1253), 
        .B2(\RegFilePlugin_regFile[7][11] ), .ZN(n707) );
  aoi22d1 U1593 ( .A1(n658), .A2(\RegFilePlugin_regFile[10][11] ), .B1(n1116), 
        .B2(\RegFilePlugin_regFile[15][11] ), .ZN(n706) );
  aoi22d1 U1594 ( .A1(n1099), .A2(\RegFilePlugin_regFile[17][11] ), .B1(n779), 
        .B2(\RegFilePlugin_regFile[23][11] ), .ZN(n705) );
  aoi22d1 U1595 ( .A1(n889), .A2(\RegFilePlugin_regFile[20][11] ), .B1(n1011), 
        .B2(\RegFilePlugin_regFile[31][11] ), .ZN(n704) );
  aoi22d1 U1596 ( .A1(n1148), .A2(\RegFilePlugin_regFile[25][11] ), .B1(n1250), 
        .B2(\RegFilePlugin_regFile[6][11] ), .ZN(n711) );
  aoi22d1 U1597 ( .A1(n1094), .A2(\RegFilePlugin_regFile[29][11] ), .B1(n1272), 
        .B2(\RegFilePlugin_regFile[11][11] ), .ZN(n710) );
  aoi22d1 U1598 ( .A1(n1073), .A2(\RegFilePlugin_regFile[2][11] ), .B1(n841), 
        .B2(\RegFilePlugin_regFile[9][11] ), .ZN(n709) );
  aoi22d1 U1599 ( .A1(n757), .A2(\RegFilePlugin_regFile[5][11] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][11] ), .ZN(n708) );
  or04d0 U1600 ( .A1(n715), .A2(n714), .A3(n713), .A4(n712), .Z(N843) );
  aoi22d1 U1601 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][2] ), .B1(n1294), 
        .B2(\RegFilePlugin_regFile[8][2] ), .ZN(n719) );
  aoi22d1 U1602 ( .A1(n1166), .A2(\RegFilePlugin_regFile[5][2] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][2] ), .ZN(n718) );
  aoi22d1 U1603 ( .A1(n1288), .A2(\RegFilePlugin_regFile[22][2] ), .B1(n1094), 
        .B2(\RegFilePlugin_regFile[29][2] ), .ZN(n717) );
  aoi22d1 U1604 ( .A1(n889), .A2(\RegFilePlugin_regFile[20][2] ), .B1(n1250), 
        .B2(\RegFilePlugin_regFile[6][2] ), .ZN(n716) );
  aoi22d1 U1605 ( .A1(n1138), .A2(\RegFilePlugin_regFile[26][2] ), .B1(n1176), 
        .B2(\RegFilePlugin_regFile[2][2] ), .ZN(n723) );
  aoi22d1 U1606 ( .A1(n1208), .A2(\RegFilePlugin_regFile[10][2] ), .B1(n926), 
        .B2(\RegFilePlugin_regFile[0][2] ), .ZN(n722) );
  aoi22d1 U1607 ( .A1(n1072), .A2(\RegFilePlugin_regFile[13][2] ), .B1(n1258), 
        .B2(\RegFilePlugin_regFile[21][2] ), .ZN(n721) );
  aoi22d1 U1608 ( .A1(n1190), .A2(\RegFilePlugin_regFile[19][2] ), .B1(n1259), 
        .B2(\RegFilePlugin_regFile[1][2] ), .ZN(n720) );
  aoi22d1 U1609 ( .A1(n884), .A2(\RegFilePlugin_regFile[12][2] ), .B1(n1011), 
        .B2(\RegFilePlugin_regFile[31][2] ), .ZN(n727) );
  aoi22d1 U1610 ( .A1(n1289), .A2(\RegFilePlugin_regFile[7][2] ), .B1(n1229), 
        .B2(\RegFilePlugin_regFile[9][2] ), .ZN(n726) );
  aoi22d1 U1611 ( .A1(n1148), .A2(\RegFilePlugin_regFile[25][2] ), .B1(n1270), 
        .B2(\RegFilePlugin_regFile[27][2] ), .ZN(n725) );
  aoi22d1 U1612 ( .A1(n1209), .A2(\RegFilePlugin_regFile[15][2] ), .B1(n1171), 
        .B2(\RegFilePlugin_regFile[11][2] ), .ZN(n724) );
  aoi22d1 U1613 ( .A1(n867), .A2(\RegFilePlugin_regFile[24][2] ), .B1(n779), 
        .B2(\RegFilePlugin_regFile[23][2] ), .ZN(n731) );
  aoi22d1 U1614 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][2] ), .B1(n1280), 
        .B2(\RegFilePlugin_regFile[3][2] ), .ZN(n730) );
  aoi22d1 U1615 ( .A1(n1217), .A2(\RegFilePlugin_regFile[4][2] ), .B1(n988), 
        .B2(\RegFilePlugin_regFile[28][2] ), .ZN(n729) );
  aoi22d1 U1616 ( .A1(n653), .A2(\RegFilePlugin_regFile[30][2] ), .B1(n1297), 
        .B2(\RegFilePlugin_regFile[18][2] ), .ZN(n728) );
  or04d0 U1617 ( .A1(n735), .A2(n734), .A3(n733), .A4(n732), .Z(N852) );
  aoi22d1 U1618 ( .A1(n1209), .A2(\RegFilePlugin_regFile[15][29] ), .B1(n1296), 
        .B2(\RegFilePlugin_regFile[12][29] ), .ZN(n740) );
  aoi22d1 U1619 ( .A1(n1244), .A2(\RegFilePlugin_regFile[13][29] ), .B1(n842), 
        .B2(\RegFilePlugin_regFile[25][29] ), .ZN(n739) );
  aoi22d1 U1620 ( .A1(n736), .A2(\RegFilePlugin_regFile[14][29] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][29] ), .ZN(n738) );
  aoi22d1 U1621 ( .A1(n1252), .A2(\RegFilePlugin_regFile[27][29] ), .B1(n1010), 
        .B2(\RegFilePlugin_regFile[16][29] ), .ZN(n737) );
  aoi22d1 U1622 ( .A1(n1288), .A2(\RegFilePlugin_regFile[22][29] ), .B1(n841), 
        .B2(\RegFilePlugin_regFile[9][29] ), .ZN(n744) );
  aoi22d1 U1623 ( .A1(n1253), .A2(\RegFilePlugin_regFile[7][29] ), .B1(n757), 
        .B2(\RegFilePlugin_regFile[5][29] ), .ZN(n743) );
  aoi22d1 U1624 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][29] ), .B1(n1258), 
        .B2(\RegFilePlugin_regFile[21][29] ), .ZN(n742) );
  aoi22d1 U1625 ( .A1(n1280), .A2(\RegFilePlugin_regFile[3][29] ), .B1(n867), 
        .B2(\RegFilePlugin_regFile[24][29] ), .ZN(n741) );
  aoi22d1 U1626 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][29] ), .B1(n1238), 
        .B2(\RegFilePlugin_regFile[4][29] ), .ZN(n748) );
  aoi22d1 U1627 ( .A1(n1269), .A2(\RegFilePlugin_regFile[1][29] ), .B1(n653), 
        .B2(\RegFilePlugin_regFile[30][29] ), .ZN(n747) );
  aoi22d1 U1628 ( .A1(n1208), .A2(\RegFilePlugin_regFile[10][29] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][29] ), .ZN(n746) );
  aoi22d1 U1629 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][29] ), .B1(n988), 
        .B2(\RegFilePlugin_regFile[28][29] ), .ZN(n745) );
  aoi22d1 U1630 ( .A1(n1222), .A2(\RegFilePlugin_regFile[20][29] ), .B1(n1176), 
        .B2(\RegFilePlugin_regFile[2][29] ), .ZN(n752) );
  aoi22d1 U1631 ( .A1(n1094), .A2(\RegFilePlugin_regFile[29][29] ), .B1(n1275), 
        .B2(\RegFilePlugin_regFile[6][29] ), .ZN(n751) );
  aoi22d1 U1632 ( .A1(n926), .A2(\RegFilePlugin_regFile[0][29] ), .B1(n1281), 
        .B2(\RegFilePlugin_regFile[23][29] ), .ZN(n750) );
  aoi22d1 U1633 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][29] ), .B1(n1171), 
        .B2(\RegFilePlugin_regFile[11][29] ), .ZN(n749) );
  or04d0 U1634 ( .A1(n756), .A2(n755), .A3(n754), .A4(n753), .Z(N825) );
  aoi22d1 U1635 ( .A1(n1210), .A2(\RegFilePlugin_regFile[3][1] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][1] ), .ZN(n762) );
  aoi22d1 U1636 ( .A1(n653), .A2(\RegFilePlugin_regFile[30][1] ), .B1(n757), 
        .B2(\RegFilePlugin_regFile[5][1] ), .ZN(n761) );
  aoi22d1 U1637 ( .A1(n758), .A2(\RegFilePlugin_regFile[19][1] ), .B1(n779), 
        .B2(\RegFilePlugin_regFile[23][1] ), .ZN(n760) );
  aoi22d1 U1638 ( .A1(n1271), .A2(\RegFilePlugin_regFile[29][1] ), .B1(n1296), 
        .B2(\RegFilePlugin_regFile[12][1] ), .ZN(n759) );
  aoi22d1 U1639 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][1] ), .B1(n988), 
        .B2(\RegFilePlugin_regFile[28][1] ), .ZN(n766) );
  aoi22d1 U1640 ( .A1(n1238), .A2(\RegFilePlugin_regFile[4][1] ), .B1(n1252), 
        .B2(\RegFilePlugin_regFile[27][1] ), .ZN(n765) );
  aoi22d1 U1641 ( .A1(n1176), .A2(\RegFilePlugin_regFile[2][1] ), .B1(n1143), 
        .B2(\RegFilePlugin_regFile[22][1] ), .ZN(n764) );
  aoi22d1 U1642 ( .A1(n1244), .A2(\RegFilePlugin_regFile[13][1] ), .B1(n1011), 
        .B2(\RegFilePlugin_regFile[31][1] ), .ZN(n763) );
  aoi22d1 U1643 ( .A1(n1253), .A2(\RegFilePlugin_regFile[7][1] ), .B1(n1295), 
        .B2(\RegFilePlugin_regFile[21][1] ), .ZN(n770) );
  aoi22d1 U1644 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][1] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][1] ), .ZN(n769) );
  aoi22d1 U1645 ( .A1(n1148), .A2(\RegFilePlugin_regFile[25][1] ), .B1(n1229), 
        .B2(\RegFilePlugin_regFile[9][1] ), .ZN(n768) );
  aoi22d1 U1646 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][1] ), .B1(n1272), 
        .B2(\RegFilePlugin_regFile[11][1] ), .ZN(n767) );
  aoi22d1 U1647 ( .A1(n1250), .A2(\RegFilePlugin_regFile[6][1] ), .B1(n1209), 
        .B2(\RegFilePlugin_regFile[15][1] ), .ZN(n774) );
  aoi22d1 U1648 ( .A1(n1273), .A2(\RegFilePlugin_regFile[24][1] ), .B1(n926), 
        .B2(\RegFilePlugin_regFile[0][1] ), .ZN(n773) );
  aoi22d1 U1649 ( .A1(n1294), .A2(\RegFilePlugin_regFile[8][1] ), .B1(n1208), 
        .B2(\RegFilePlugin_regFile[10][1] ), .ZN(n772) );
  aoi22d1 U1650 ( .A1(n889), .A2(\RegFilePlugin_regFile[20][1] ), .B1(n1259), 
        .B2(\RegFilePlugin_regFile[1][1] ), .ZN(n771) );
  or04d0 U1651 ( .A1(n778), .A2(n777), .A3(n776), .A4(n775), .Z(N853) );
  aoi22d1 U1652 ( .A1(n1116), .A2(\RegFilePlugin_regFile[15][17] ), .B1(n1295), 
        .B2(\RegFilePlugin_regFile[21][17] ), .ZN(n784) );
  aoi22d1 U1653 ( .A1(n1148), .A2(\RegFilePlugin_regFile[25][17] ), .B1(n779), 
        .B2(\RegFilePlugin_regFile[23][17] ), .ZN(n783) );
  aoi22d1 U1654 ( .A1(n1289), .A2(\RegFilePlugin_regFile[7][17] ), .B1(n780), 
        .B2(\RegFilePlugin_regFile[27][17] ), .ZN(n782) );
  aoi22d1 U1655 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][17] ), .B1(n1260), 
        .B2(\RegFilePlugin_regFile[30][17] ), .ZN(n781) );
  aoi22d1 U1656 ( .A1(n1238), .A2(\RegFilePlugin_regFile[4][17] ), .B1(n1296), 
        .B2(\RegFilePlugin_regFile[12][17] ), .ZN(n788) );
  aoi22d1 U1657 ( .A1(n1273), .A2(\RegFilePlugin_regFile[24][17] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][17] ), .ZN(n787) );
  aoi22d1 U1658 ( .A1(n1099), .A2(\RegFilePlugin_regFile[17][17] ), .B1(n1272), 
        .B2(\RegFilePlugin_regFile[11][17] ), .ZN(n786) );
  aoi22d1 U1659 ( .A1(n1298), .A2(\RegFilePlugin_regFile[28][17] ), .B1(n841), 
        .B2(\RegFilePlugin_regFile[9][17] ), .ZN(n785) );
  aoi22d1 U1660 ( .A1(n1244), .A2(\RegFilePlugin_regFile[13][17] ), .B1(n1222), 
        .B2(\RegFilePlugin_regFile[20][17] ), .ZN(n792) );
  aoi22d1 U1661 ( .A1(n1094), .A2(\RegFilePlugin_regFile[29][17] ), .B1(n926), 
        .B2(\RegFilePlugin_regFile[0][17] ), .ZN(n791) );
  aoi22d1 U1662 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][17] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][17] ), .ZN(n790) );
  aoi22d1 U1663 ( .A1(n1275), .A2(\RegFilePlugin_regFile[6][17] ), .B1(n1011), 
        .B2(\RegFilePlugin_regFile[31][17] ), .ZN(n789) );
  aoi22d1 U1664 ( .A1(n1073), .A2(\RegFilePlugin_regFile[2][17] ), .B1(n757), 
        .B2(\RegFilePlugin_regFile[5][17] ), .ZN(n796) );
  aoi22d1 U1665 ( .A1(n1143), .A2(\RegFilePlugin_regFile[22][17] ), .B1(n1210), 
        .B2(\RegFilePlugin_regFile[3][17] ), .ZN(n795) );
  aoi22d1 U1666 ( .A1(n1294), .A2(\RegFilePlugin_regFile[8][17] ), .B1(n1269), 
        .B2(\RegFilePlugin_regFile[1][17] ), .ZN(n794) );
  aoi22d1 U1667 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][17] ), .B1(n658), 
        .B2(\RegFilePlugin_regFile[10][17] ), .ZN(n793) );
  or04d0 U1668 ( .A1(n800), .A2(n799), .A3(n798), .A4(n797), .Z(N837) );
  aoi22d1 U1669 ( .A1(n1280), .A2(\RegFilePlugin_regFile[3][22] ), .B1(n1272), 
        .B2(\RegFilePlugin_regFile[11][22] ), .ZN(n804) );
  aoi22d1 U1670 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][22] ), .B1(n1148), 
        .B2(\RegFilePlugin_regFile[25][22] ), .ZN(n803) );
  aoi22d1 U1671 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][22] ), .B1(n1298), 
        .B2(\RegFilePlugin_regFile[28][22] ), .ZN(n802) );
  aoi22d1 U1672 ( .A1(n1176), .A2(\RegFilePlugin_regFile[2][22] ), .B1(n1011), 
        .B2(\RegFilePlugin_regFile[31][22] ), .ZN(n801) );
  aoi22d1 U1673 ( .A1(n1094), .A2(\RegFilePlugin_regFile[29][22] ), .B1(n1258), 
        .B2(\RegFilePlugin_regFile[21][22] ), .ZN(n808) );
  aoi22d1 U1674 ( .A1(n1099), .A2(\RegFilePlugin_regFile[17][22] ), .B1(n1273), 
        .B2(\RegFilePlugin_regFile[24][22] ), .ZN(n807) );
  aoi22d1 U1675 ( .A1(n1259), .A2(\RegFilePlugin_regFile[1][22] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][22] ), .ZN(n806) );
  aoi22d1 U1676 ( .A1(n757), .A2(\RegFilePlugin_regFile[5][22] ), .B1(n1217), 
        .B2(\RegFilePlugin_regFile[4][22] ), .ZN(n805) );
  aoi22d1 U1677 ( .A1(n1208), .A2(\RegFilePlugin_regFile[10][22] ), .B1(n926), 
        .B2(\RegFilePlugin_regFile[0][22] ), .ZN(n812) );
  aoi22d1 U1678 ( .A1(n1072), .A2(\RegFilePlugin_regFile[13][22] ), .B1(n1252), 
        .B2(\RegFilePlugin_regFile[27][22] ), .ZN(n811) );
  aoi22d1 U1679 ( .A1(n1138), .A2(\RegFilePlugin_regFile[26][22] ), .B1(n1260), 
        .B2(\RegFilePlugin_regFile[30][22] ), .ZN(n810) );
  aoi22d1 U1680 ( .A1(n1250), .A2(\RegFilePlugin_regFile[6][22] ), .B1(n841), 
        .B2(\RegFilePlugin_regFile[9][22] ), .ZN(n809) );
  aoi22d1 U1681 ( .A1(n1209), .A2(\RegFilePlugin_regFile[15][22] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][22] ), .ZN(n816) );
  aoi22d1 U1682 ( .A1(n1222), .A2(\RegFilePlugin_regFile[20][22] ), .B1(n1282), 
        .B2(\RegFilePlugin_regFile[14][22] ), .ZN(n815) );
  aoi22d1 U1683 ( .A1(n1289), .A2(\RegFilePlugin_regFile[7][22] ), .B1(n1281), 
        .B2(\RegFilePlugin_regFile[23][22] ), .ZN(n814) );
  aoi22d1 U1684 ( .A1(n1143), .A2(\RegFilePlugin_regFile[22][22] ), .B1(n884), 
        .B2(\RegFilePlugin_regFile[12][22] ), .ZN(n813) );
  or04d0 U1685 ( .A1(n820), .A2(n819), .A3(n818), .A4(n817), .Z(N832) );
  aoi22d1 U1686 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][6] ), .B1(n1272), 
        .B2(\RegFilePlugin_regFile[11][6] ), .ZN(n824) );
  aoi22d1 U1687 ( .A1(n1148), .A2(\RegFilePlugin_regFile[25][6] ), .B1(n1116), 
        .B2(\RegFilePlugin_regFile[15][6] ), .ZN(n823) );
  aoi22d1 U1688 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][6] ), .B1(n1269), 
        .B2(\RegFilePlugin_regFile[1][6] ), .ZN(n822) );
  aoi22d1 U1689 ( .A1(n1094), .A2(\RegFilePlugin_regFile[29][6] ), .B1(n1010), 
        .B2(\RegFilePlugin_regFile[16][6] ), .ZN(n821) );
  aoi22d1 U1690 ( .A1(n658), .A2(\RegFilePlugin_regFile[10][6] ), .B1(n926), 
        .B2(\RegFilePlugin_regFile[0][6] ), .ZN(n828) );
  aoi22d1 U1691 ( .A1(n653), .A2(\RegFilePlugin_regFile[30][6] ), .B1(n1297), 
        .B2(\RegFilePlugin_regFile[18][6] ), .ZN(n827) );
  aoi22d1 U1692 ( .A1(n1294), .A2(\RegFilePlugin_regFile[8][6] ), .B1(n1298), 
        .B2(\RegFilePlugin_regFile[28][6] ), .ZN(n826) );
  aoi22d1 U1693 ( .A1(n1222), .A2(\RegFilePlugin_regFile[20][6] ), .B1(n779), 
        .B2(\RegFilePlugin_regFile[23][6] ), .ZN(n825) );
  aoi22d1 U1694 ( .A1(n1217), .A2(\RegFilePlugin_regFile[4][6] ), .B1(n1295), 
        .B2(\RegFilePlugin_regFile[21][6] ), .ZN(n832) );
  aoi22d1 U1695 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][6] ), .B1(n1143), 
        .B2(\RegFilePlugin_regFile[22][6] ), .ZN(n831) );
  aoi22d1 U1696 ( .A1(n1073), .A2(\RegFilePlugin_regFile[2][6] ), .B1(n841), 
        .B2(\RegFilePlugin_regFile[9][6] ), .ZN(n830) );
  aoi22d1 U1697 ( .A1(n1244), .A2(\RegFilePlugin_regFile[13][6] ), .B1(n884), 
        .B2(\RegFilePlugin_regFile[12][6] ), .ZN(n829) );
  aoi22d1 U1698 ( .A1(n1190), .A2(\RegFilePlugin_regFile[19][6] ), .B1(n1270), 
        .B2(\RegFilePlugin_regFile[27][6] ), .ZN(n836) );
  aoi22d1 U1699 ( .A1(n1253), .A2(\RegFilePlugin_regFile[7][6] ), .B1(n1166), 
        .B2(\RegFilePlugin_regFile[5][6] ), .ZN(n835) );
  aoi22d1 U1700 ( .A1(n1275), .A2(\RegFilePlugin_regFile[6][6] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][6] ), .ZN(n834) );
  aoi22d1 U1701 ( .A1(n1280), .A2(\RegFilePlugin_regFile[3][6] ), .B1(n1273), 
        .B2(\RegFilePlugin_regFile[24][6] ), .ZN(n833) );
  or04d0 U1702 ( .A1(n840), .A2(n839), .A3(n838), .A4(n837), .Z(N848) );
  aoi22d1 U1703 ( .A1(n1271), .A2(\RegFilePlugin_regFile[29][13] ), .B1(n841), 
        .B2(\RegFilePlugin_regFile[9][13] ), .ZN(n846) );
  aoi22d1 U1704 ( .A1(n842), .A2(\RegFilePlugin_regFile[25][13] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][13] ), .ZN(n845) );
  aoi22d1 U1705 ( .A1(n1250), .A2(\RegFilePlugin_regFile[6][13] ), .B1(n884), 
        .B2(\RegFilePlugin_regFile[12][13] ), .ZN(n844) );
  aoi22d1 U1706 ( .A1(n1072), .A2(\RegFilePlugin_regFile[13][13] ), .B1(n1295), 
        .B2(\RegFilePlugin_regFile[21][13] ), .ZN(n843) );
  aoi22d1 U1707 ( .A1(n1166), .A2(\RegFilePlugin_regFile[5][13] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][13] ), .ZN(n850) );
  aoi22d1 U1708 ( .A1(n1073), .A2(\RegFilePlugin_regFile[2][13] ), .B1(n1210), 
        .B2(\RegFilePlugin_regFile[3][13] ), .ZN(n849) );
  aoi22d1 U1709 ( .A1(n889), .A2(\RegFilePlugin_regFile[20][13] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][13] ), .ZN(n848) );
  aoi22d1 U1710 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][13] ), .B1(n1209), 
        .B2(\RegFilePlugin_regFile[15][13] ), .ZN(n847) );
  aoi22d1 U1711 ( .A1(n658), .A2(\RegFilePlugin_regFile[10][13] ), .B1(n988), 
        .B2(\RegFilePlugin_regFile[28][13] ), .ZN(n854) );
  aoi22d1 U1712 ( .A1(n1294), .A2(\RegFilePlugin_regFile[8][13] ), .B1(n1269), 
        .B2(\RegFilePlugin_regFile[1][13] ), .ZN(n853) );
  aoi22d1 U1713 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][13] ), .B1(n779), 
        .B2(\RegFilePlugin_regFile[23][13] ), .ZN(n852) );
  aoi22d1 U1714 ( .A1(n1273), .A2(\RegFilePlugin_regFile[24][13] ), .B1(n1252), 
        .B2(\RegFilePlugin_regFile[27][13] ), .ZN(n851) );
  aoi22d1 U1715 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][13] ), .B1(n1272), 
        .B2(\RegFilePlugin_regFile[11][13] ), .ZN(n858) );
  aoi22d1 U1716 ( .A1(n1288), .A2(\RegFilePlugin_regFile[22][13] ), .B1(n653), 
        .B2(\RegFilePlugin_regFile[30][13] ), .ZN(n857) );
  aoi22d1 U1717 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][13] ), .B1(n1217), 
        .B2(\RegFilePlugin_regFile[4][13] ), .ZN(n856) );
  aoi22d1 U1718 ( .A1(n1289), .A2(\RegFilePlugin_regFile[7][13] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][13] ), .ZN(n855) );
  or04d0 U1719 ( .A1(n862), .A2(n861), .A3(n860), .A4(n859), .Z(N841) );
  aoi22d1 U1720 ( .A1(n1073), .A2(\RegFilePlugin_regFile[2][20] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][20] ), .ZN(n866) );
  aoi22d1 U1721 ( .A1(n1282), .A2(\RegFilePlugin_regFile[14][20] ), .B1(n1289), 
        .B2(\RegFilePlugin_regFile[7][20] ), .ZN(n865) );
  aoi22d1 U1722 ( .A1(n1138), .A2(\RegFilePlugin_regFile[26][20] ), .B1(n1148), 
        .B2(\RegFilePlugin_regFile[25][20] ), .ZN(n864) );
  aoi22d1 U1723 ( .A1(n1298), .A2(\RegFilePlugin_regFile[28][20] ), .B1(n1281), 
        .B2(\RegFilePlugin_regFile[23][20] ), .ZN(n863) );
  aoi22d1 U1724 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][20] ), .B1(n1269), 
        .B2(\RegFilePlugin_regFile[1][20] ), .ZN(n871) );
  aoi22d1 U1725 ( .A1(n867), .A2(\RegFilePlugin_regFile[24][20] ), .B1(n1252), 
        .B2(\RegFilePlugin_regFile[27][20] ), .ZN(n870) );
  aoi22d1 U1726 ( .A1(n926), .A2(\RegFilePlugin_regFile[0][20] ), .B1(n1229), 
        .B2(\RegFilePlugin_regFile[9][20] ), .ZN(n869) );
  aoi22d1 U1727 ( .A1(n1250), .A2(\RegFilePlugin_regFile[6][20] ), .B1(n1296), 
        .B2(\RegFilePlugin_regFile[12][20] ), .ZN(n868) );
  aoi22d1 U1728 ( .A1(n1072), .A2(\RegFilePlugin_regFile[13][20] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][20] ), .ZN(n875) );
  aoi22d1 U1729 ( .A1(n1260), .A2(\RegFilePlugin_regFile[30][20] ), .B1(n1295), 
        .B2(\RegFilePlugin_regFile[21][20] ), .ZN(n874) );
  aoi22d1 U1730 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][20] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][20] ), .ZN(n873) );
  aoi22d1 U1731 ( .A1(n889), .A2(\RegFilePlugin_regFile[20][20] ), .B1(n1143), 
        .B2(\RegFilePlugin_regFile[22][20] ), .ZN(n872) );
  aoi22d1 U1732 ( .A1(n1094), .A2(\RegFilePlugin_regFile[29][20] ), .B1(n1209), 
        .B2(\RegFilePlugin_regFile[15][20] ), .ZN(n879) );
  aoi22d1 U1733 ( .A1(n1099), .A2(\RegFilePlugin_regFile[17][20] ), .B1(n1217), 
        .B2(\RegFilePlugin_regFile[4][20] ), .ZN(n878) );
  aoi22d1 U1734 ( .A1(n1280), .A2(\RegFilePlugin_regFile[3][20] ), .B1(n1171), 
        .B2(\RegFilePlugin_regFile[11][20] ), .ZN(n877) );
  aoi22d1 U1735 ( .A1(n658), .A2(\RegFilePlugin_regFile[10][20] ), .B1(n757), 
        .B2(\RegFilePlugin_regFile[5][20] ), .ZN(n876) );
  or04d0 U1736 ( .A1(n883), .A2(n882), .A3(n881), .A4(n880), .Z(N834) );
  aoi22d1 U1737 ( .A1(n1116), .A2(\RegFilePlugin_regFile[15][24] ), .B1(n884), 
        .B2(\RegFilePlugin_regFile[12][24] ), .ZN(n888) );
  aoi22d1 U1738 ( .A1(n1297), .A2(\RegFilePlugin_regFile[18][24] ), .B1(n1229), 
        .B2(\RegFilePlugin_regFile[9][24] ), .ZN(n887) );
  aoi22d1 U1739 ( .A1(n1148), .A2(\RegFilePlugin_regFile[25][24] ), .B1(n1289), 
        .B2(\RegFilePlugin_regFile[7][24] ), .ZN(n886) );
  aoi22d1 U1740 ( .A1(n1190), .A2(\RegFilePlugin_regFile[19][24] ), .B1(n1273), 
        .B2(\RegFilePlugin_regFile[24][24] ), .ZN(n885) );
  aoi22d1 U1741 ( .A1(n1288), .A2(\RegFilePlugin_regFile[22][24] ), .B1(n1217), 
        .B2(\RegFilePlugin_regFile[4][24] ), .ZN(n893) );
  aoi22d1 U1742 ( .A1(n1208), .A2(\RegFilePlugin_regFile[10][24] ), .B1(n1280), 
        .B2(\RegFilePlugin_regFile[3][24] ), .ZN(n892) );
  aoi22d1 U1743 ( .A1(n889), .A2(\RegFilePlugin_regFile[20][24] ), .B1(n1281), 
        .B2(\RegFilePlugin_regFile[23][24] ), .ZN(n891) );
  aoi22d1 U1744 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][24] ), .B1(n1171), 
        .B2(\RegFilePlugin_regFile[11][24] ), .ZN(n890) );
  aoi22d1 U1745 ( .A1(n1275), .A2(\RegFilePlugin_regFile[6][24] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][24] ), .ZN(n897) );
  aoi22d1 U1746 ( .A1(n1176), .A2(\RegFilePlugin_regFile[2][24] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][24] ), .ZN(n896) );
  aoi22d1 U1747 ( .A1(n1260), .A2(\RegFilePlugin_regFile[30][24] ), .B1(n988), 
        .B2(\RegFilePlugin_regFile[28][24] ), .ZN(n895) );
  aoi22d1 U1748 ( .A1(n1166), .A2(\RegFilePlugin_regFile[5][24] ), .B1(n1258), 
        .B2(\RegFilePlugin_regFile[21][24] ), .ZN(n894) );
  aoi22d1 U1749 ( .A1(n1282), .A2(\RegFilePlugin_regFile[14][24] ), .B1(n1269), 
        .B2(\RegFilePlugin_regFile[1][24] ), .ZN(n901) );
  aoi22d1 U1750 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][24] ), .B1(n1252), 
        .B2(\RegFilePlugin_regFile[27][24] ), .ZN(n900) );
  aoi22d1 U1751 ( .A1(n1271), .A2(\RegFilePlugin_regFile[29][24] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][24] ), .ZN(n899) );
  aoi22d1 U1752 ( .A1(n1138), .A2(\RegFilePlugin_regFile[26][24] ), .B1(n1244), 
        .B2(\RegFilePlugin_regFile[13][24] ), .ZN(n898) );
  or04d0 U1753 ( .A1(n905), .A2(n904), .A3(n903), .A4(n902), .Z(N830) );
  aoi22d1 U1754 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][5] ), .B1(n1271), 
        .B2(\RegFilePlugin_regFile[29][5] ), .ZN(n909) );
  aoi22d1 U1755 ( .A1(n1143), .A2(\RegFilePlugin_regFile[22][5] ), .B1(n779), 
        .B2(\RegFilePlugin_regFile[23][5] ), .ZN(n908) );
  aoi22d1 U1756 ( .A1(n1238), .A2(\RegFilePlugin_regFile[4][5] ), .B1(n1250), 
        .B2(\RegFilePlugin_regFile[6][5] ), .ZN(n907) );
  aoi22d1 U1757 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][5] ), .B1(n926), 
        .B2(\RegFilePlugin_regFile[0][5] ), .ZN(n906) );
  aoi22d1 U1758 ( .A1(n1269), .A2(\RegFilePlugin_regFile[1][5] ), .B1(n653), 
        .B2(\RegFilePlugin_regFile[30][5] ), .ZN(n913) );
  aoi22d1 U1759 ( .A1(n889), .A2(\RegFilePlugin_regFile[20][5] ), .B1(n884), 
        .B2(\RegFilePlugin_regFile[12][5] ), .ZN(n912) );
  aoi22d1 U1760 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][5] ), .B1(n1270), 
        .B2(\RegFilePlugin_regFile[27][5] ), .ZN(n911) );
  aoi22d1 U1761 ( .A1(n658), .A2(\RegFilePlugin_regFile[10][5] ), .B1(n988), 
        .B2(\RegFilePlugin_regFile[28][5] ), .ZN(n910) );
  aoi22d1 U1762 ( .A1(n1190), .A2(\RegFilePlugin_regFile[19][5] ), .B1(n1229), 
        .B2(\RegFilePlugin_regFile[9][5] ), .ZN(n917) );
  aoi22d1 U1763 ( .A1(n1116), .A2(\RegFilePlugin_regFile[15][5] ), .B1(n1010), 
        .B2(\RegFilePlugin_regFile[16][5] ), .ZN(n916) );
  aoi22d1 U1764 ( .A1(n1280), .A2(\RegFilePlugin_regFile[3][5] ), .B1(n1295), 
        .B2(\RegFilePlugin_regFile[21][5] ), .ZN(n915) );
  aoi22d1 U1765 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][5] ), .B1(n867), 
        .B2(\RegFilePlugin_regFile[24][5] ), .ZN(n914) );
  aoi22d1 U1766 ( .A1(n1073), .A2(\RegFilePlugin_regFile[2][5] ), .B1(n1272), 
        .B2(\RegFilePlugin_regFile[11][5] ), .ZN(n921) );
  aoi22d1 U1767 ( .A1(n1166), .A2(\RegFilePlugin_regFile[5][5] ), .B1(n1011), 
        .B2(\RegFilePlugin_regFile[31][5] ), .ZN(n920) );
  aoi22d1 U1768 ( .A1(n1244), .A2(\RegFilePlugin_regFile[13][5] ), .B1(n1297), 
        .B2(\RegFilePlugin_regFile[18][5] ), .ZN(n919) );
  aoi22d1 U1769 ( .A1(n1148), .A2(\RegFilePlugin_regFile[25][5] ), .B1(n1253), 
        .B2(\RegFilePlugin_regFile[7][5] ), .ZN(n918) );
  or04d0 U1770 ( .A1(n925), .A2(n924), .A3(n923), .A4(n922), .Z(N849) );
  aoi22d1 U1771 ( .A1(n926), .A2(\RegFilePlugin_regFile[0][3] ), .B1(n779), 
        .B2(\RegFilePlugin_regFile[23][3] ), .ZN(n930) );
  aoi22d1 U1772 ( .A1(n1298), .A2(\RegFilePlugin_regFile[28][3] ), .B1(n1011), 
        .B2(\RegFilePlugin_regFile[31][3] ), .ZN(n929) );
  aoi22d1 U1773 ( .A1(n1138), .A2(\RegFilePlugin_regFile[26][3] ), .B1(n1270), 
        .B2(\RegFilePlugin_regFile[27][3] ), .ZN(n928) );
  aoi22d1 U1774 ( .A1(n1244), .A2(\RegFilePlugin_regFile[13][3] ), .B1(n1294), 
        .B2(\RegFilePlugin_regFile[8][3] ), .ZN(n927) );
  aoi22d1 U1775 ( .A1(n1259), .A2(\RegFilePlugin_regFile[1][3] ), .B1(n1166), 
        .B2(\RegFilePlugin_regFile[5][3] ), .ZN(n934) );
  aoi22d1 U1776 ( .A1(n1099), .A2(\RegFilePlugin_regFile[17][3] ), .B1(n1208), 
        .B2(\RegFilePlugin_regFile[10][3] ), .ZN(n933) );
  aoi22d1 U1777 ( .A1(n889), .A2(\RegFilePlugin_regFile[20][3] ), .B1(n1229), 
        .B2(\RegFilePlugin_regFile[9][3] ), .ZN(n932) );
  aoi22d1 U1778 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][3] ), .B1(n842), 
        .B2(\RegFilePlugin_regFile[25][3] ), .ZN(n931) );
  aoi22d1 U1779 ( .A1(n1288), .A2(\RegFilePlugin_regFile[22][3] ), .B1(n1280), 
        .B2(\RegFilePlugin_regFile[3][3] ), .ZN(n938) );
  aoi22d1 U1780 ( .A1(n1217), .A2(\RegFilePlugin_regFile[4][3] ), .B1(n1275), 
        .B2(\RegFilePlugin_regFile[6][3] ), .ZN(n937) );
  aoi22d1 U1781 ( .A1(n867), .A2(\RegFilePlugin_regFile[24][3] ), .B1(n1295), 
        .B2(\RegFilePlugin_regFile[21][3] ), .ZN(n936) );
  aoi22d1 U1782 ( .A1(n1094), .A2(\RegFilePlugin_regFile[29][3] ), .B1(n1171), 
        .B2(\RegFilePlugin_regFile[11][3] ), .ZN(n935) );
  aoi22d1 U1783 ( .A1(n1176), .A2(\RegFilePlugin_regFile[2][3] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][3] ), .ZN(n942) );
  aoi22d1 U1784 ( .A1(n1297), .A2(\RegFilePlugin_regFile[18][3] ), .B1(n1296), 
        .B2(\RegFilePlugin_regFile[12][3] ), .ZN(n941) );
  aoi22d1 U1785 ( .A1(n1260), .A2(\RegFilePlugin_regFile[30][3] ), .B1(n1209), 
        .B2(\RegFilePlugin_regFile[15][3] ), .ZN(n940) );
  aoi22d1 U1786 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][3] ), .B1(n1253), 
        .B2(\RegFilePlugin_regFile[7][3] ), .ZN(n939) );
  or04d0 U1787 ( .A1(n946), .A2(n945), .A3(n944), .A4(n943), .Z(N851) );
  aoi22d1 U1788 ( .A1(n842), .A2(\RegFilePlugin_regFile[25][19] ), .B1(n653), 
        .B2(\RegFilePlugin_regFile[30][19] ), .ZN(n950) );
  aoi22d1 U1789 ( .A1(n1269), .A2(\RegFilePlugin_regFile[1][19] ), .B1(n884), 
        .B2(\RegFilePlugin_regFile[12][19] ), .ZN(n949) );
  aoi22d1 U1790 ( .A1(n1072), .A2(\RegFilePlugin_regFile[13][19] ), .B1(n1171), 
        .B2(\RegFilePlugin_regFile[11][19] ), .ZN(n948) );
  aoi22d1 U1791 ( .A1(n1073), .A2(\RegFilePlugin_regFile[2][19] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][19] ), .ZN(n947) );
  aoi22d1 U1792 ( .A1(n1297), .A2(\RegFilePlugin_regFile[18][19] ), .B1(n926), 
        .B2(\RegFilePlugin_regFile[0][19] ), .ZN(n954) );
  aoi22d1 U1793 ( .A1(n757), .A2(\RegFilePlugin_regFile[5][19] ), .B1(n1270), 
        .B2(\RegFilePlugin_regFile[27][19] ), .ZN(n953) );
  aoi22d1 U1794 ( .A1(n1210), .A2(\RegFilePlugin_regFile[3][19] ), .B1(n1116), 
        .B2(\RegFilePlugin_regFile[15][19] ), .ZN(n952) );
  aoi22d1 U1795 ( .A1(n1282), .A2(\RegFilePlugin_regFile[14][19] ), .B1(n1281), 
        .B2(\RegFilePlugin_regFile[23][19] ), .ZN(n951) );
  aoi22d1 U1796 ( .A1(n1143), .A2(\RegFilePlugin_regFile[22][19] ), .B1(n1229), 
        .B2(\RegFilePlugin_regFile[9][19] ), .ZN(n958) );
  aoi22d1 U1797 ( .A1(n889), .A2(\RegFilePlugin_regFile[20][19] ), .B1(n1258), 
        .B2(\RegFilePlugin_regFile[21][19] ), .ZN(n957) );
  aoi22d1 U1798 ( .A1(n1298), .A2(\RegFilePlugin_regFile[28][19] ), .B1(n867), 
        .B2(\RegFilePlugin_regFile[24][19] ), .ZN(n956) );
  aoi22d1 U1799 ( .A1(n1099), .A2(\RegFilePlugin_regFile[17][19] ), .B1(n1271), 
        .B2(\RegFilePlugin_regFile[29][19] ), .ZN(n955) );
  aoi22d1 U1800 ( .A1(n1138), .A2(\RegFilePlugin_regFile[26][19] ), .B1(n1289), 
        .B2(\RegFilePlugin_regFile[7][19] ), .ZN(n962) );
  aoi22d1 U1801 ( .A1(n658), .A2(\RegFilePlugin_regFile[10][19] ), .B1(n1238), 
        .B2(\RegFilePlugin_regFile[4][19] ), .ZN(n961) );
  aoi22d1 U1802 ( .A1(n1294), .A2(\RegFilePlugin_regFile[8][19] ), .B1(n1250), 
        .B2(\RegFilePlugin_regFile[6][19] ), .ZN(n960) );
  aoi22d1 U1803 ( .A1(n1190), .A2(\RegFilePlugin_regFile[19][19] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][19] ), .ZN(n959) );
  or04d0 U1804 ( .A1(n966), .A2(n965), .A3(n964), .A4(n963), .Z(N835) );
  aoi22d1 U1805 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][9] ), .B1(n1166), 
        .B2(\RegFilePlugin_regFile[5][9] ), .ZN(n970) );
  aoi22d1 U1806 ( .A1(n1208), .A2(\RegFilePlugin_regFile[10][9] ), .B1(n988), 
        .B2(\RegFilePlugin_regFile[28][9] ), .ZN(n969) );
  aoi22d1 U1807 ( .A1(n1073), .A2(\RegFilePlugin_regFile[2][9] ), .B1(n884), 
        .B2(\RegFilePlugin_regFile[12][9] ), .ZN(n968) );
  aoi22d1 U1808 ( .A1(n1260), .A2(\RegFilePlugin_regFile[30][9] ), .B1(n1250), 
        .B2(\RegFilePlugin_regFile[6][9] ), .ZN(n967) );
  aoi22d1 U1809 ( .A1(n889), .A2(\RegFilePlugin_regFile[20][9] ), .B1(n1238), 
        .B2(\RegFilePlugin_regFile[4][9] ), .ZN(n974) );
  aoi22d1 U1810 ( .A1(n1281), .A2(\RegFilePlugin_regFile[23][9] ), .B1(n1010), 
        .B2(\RegFilePlugin_regFile[16][9] ), .ZN(n973) );
  aoi22d1 U1811 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][9] ), .B1(n1259), 
        .B2(\RegFilePlugin_regFile[1][9] ), .ZN(n972) );
  aoi22d1 U1812 ( .A1(n1148), .A2(\RegFilePlugin_regFile[25][9] ), .B1(n867), 
        .B2(\RegFilePlugin_regFile[24][9] ), .ZN(n971) );
  aoi22d1 U1813 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][9] ), .B1(n1190), 
        .B2(\RegFilePlugin_regFile[19][9] ), .ZN(n978) );
  aoi22d1 U1814 ( .A1(n1244), .A2(\RegFilePlugin_regFile[13][9] ), .B1(n1143), 
        .B2(\RegFilePlugin_regFile[22][9] ), .ZN(n977) );
  aoi22d1 U1815 ( .A1(n1116), .A2(\RegFilePlugin_regFile[15][9] ), .B1(n1272), 
        .B2(\RegFilePlugin_regFile[11][9] ), .ZN(n976) );
  aoi22d1 U1816 ( .A1(n1094), .A2(\RegFilePlugin_regFile[29][9] ), .B1(n1270), 
        .B2(\RegFilePlugin_regFile[27][9] ), .ZN(n975) );
  aoi22d1 U1817 ( .A1(n1258), .A2(\RegFilePlugin_regFile[21][9] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][9] ), .ZN(n982) );
  aoi22d1 U1818 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][9] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][9] ), .ZN(n981) );
  aoi22d1 U1819 ( .A1(n1297), .A2(\RegFilePlugin_regFile[18][9] ), .B1(n841), 
        .B2(\RegFilePlugin_regFile[9][9] ), .ZN(n980) );
  aoi22d1 U1820 ( .A1(n1253), .A2(\RegFilePlugin_regFile[7][9] ), .B1(n1210), 
        .B2(\RegFilePlugin_regFile[3][9] ), .ZN(n979) );
  or04d0 U1821 ( .A1(n986), .A2(n985), .A3(n984), .A4(n983), .Z(N845) );
  aoi22d1 U1822 ( .A1(n1294), .A2(\RegFilePlugin_regFile[8][0] ), .B1(n779), 
        .B2(\RegFilePlugin_regFile[23][0] ), .ZN(n993) );
  aoi22d1 U1823 ( .A1(n988), .A2(\RegFilePlugin_regFile[28][0] ), .B1(n987), 
        .B2(\RegFilePlugin_regFile[21][0] ), .ZN(n992) );
  aoi22d1 U1824 ( .A1(n989), .A2(\RegFilePlugin_regFile[11][0] ), .B1(n1011), 
        .B2(\RegFilePlugin_regFile[31][0] ), .ZN(n991) );
  aoi22d1 U1825 ( .A1(n1280), .A2(\RegFilePlugin_regFile[3][0] ), .B1(n1250), 
        .B2(\RegFilePlugin_regFile[6][0] ), .ZN(n990) );
  aoi22d1 U1826 ( .A1(n1273), .A2(\RegFilePlugin_regFile[24][0] ), .B1(n1252), 
        .B2(\RegFilePlugin_regFile[27][0] ), .ZN(n997) );
  aoi22d1 U1827 ( .A1(n1143), .A2(\RegFilePlugin_regFile[22][0] ), .B1(n1297), 
        .B2(\RegFilePlugin_regFile[18][0] ), .ZN(n996) );
  aoi22d1 U1828 ( .A1(n1244), .A2(\RegFilePlugin_regFile[13][0] ), .B1(n1229), 
        .B2(\RegFilePlugin_regFile[9][0] ), .ZN(n995) );
  aoi22d1 U1829 ( .A1(n1222), .A2(\RegFilePlugin_regFile[20][0] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][0] ), .ZN(n994) );
  aoi22d1 U1830 ( .A1(n1259), .A2(\RegFilePlugin_regFile[1][0] ), .B1(n926), 
        .B2(\RegFilePlugin_regFile[0][0] ), .ZN(n1001) );
  aoi22d1 U1831 ( .A1(n1138), .A2(\RegFilePlugin_regFile[26][0] ), .B1(n1094), 
        .B2(\RegFilePlugin_regFile[29][0] ), .ZN(n1000) );
  aoi22d1 U1832 ( .A1(n1260), .A2(\RegFilePlugin_regFile[30][0] ), .B1(n884), 
        .B2(\RegFilePlugin_regFile[12][0] ), .ZN(n999) );
  aoi22d1 U1833 ( .A1(n1282), .A2(\RegFilePlugin_regFile[14][0] ), .B1(n757), 
        .B2(\RegFilePlugin_regFile[5][0] ), .ZN(n998) );
  aoi22d1 U1834 ( .A1(n658), .A2(\RegFilePlugin_regFile[10][0] ), .B1(n1238), 
        .B2(\RegFilePlugin_regFile[4][0] ), .ZN(n1005) );
  aoi22d1 U1835 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][0] ), .B1(n1116), 
        .B2(\RegFilePlugin_regFile[15][0] ), .ZN(n1004) );
  aoi22d1 U1836 ( .A1(n1190), .A2(\RegFilePlugin_regFile[19][0] ), .B1(n1253), 
        .B2(\RegFilePlugin_regFile[7][0] ), .ZN(n1003) );
  aoi22d1 U1837 ( .A1(n842), .A2(\RegFilePlugin_regFile[25][0] ), .B1(n1176), 
        .B2(\RegFilePlugin_regFile[2][0] ), .ZN(n1002) );
  or04d0 U1838 ( .A1(n1009), .A2(n1008), .A3(n1007), .A4(n1006), .Z(N854) );
  aoi22d1 U1839 ( .A1(n1094), .A2(\RegFilePlugin_regFile[29][16] ), .B1(n1010), 
        .B2(\RegFilePlugin_regFile[16][16] ), .ZN(n1015) );
  aoi22d1 U1840 ( .A1(n779), .A2(\RegFilePlugin_regFile[23][16] ), .B1(n1011), 
        .B2(\RegFilePlugin_regFile[31][16] ), .ZN(n1014) );
  aoi22d1 U1841 ( .A1(n1222), .A2(\RegFilePlugin_regFile[20][16] ), .B1(n1210), 
        .B2(\RegFilePlugin_regFile[3][16] ), .ZN(n1013) );
  aoi22d1 U1842 ( .A1(n1282), .A2(\RegFilePlugin_regFile[14][16] ), .B1(n1289), 
        .B2(\RegFilePlugin_regFile[7][16] ), .ZN(n1012) );
  aoi22d1 U1843 ( .A1(n1294), .A2(\RegFilePlugin_regFile[8][16] ), .B1(n1250), 
        .B2(\RegFilePlugin_regFile[6][16] ), .ZN(n1019) );
  aoi22d1 U1844 ( .A1(n842), .A2(\RegFilePlugin_regFile[25][16] ), .B1(n1252), 
        .B2(\RegFilePlugin_regFile[27][16] ), .ZN(n1018) );
  aoi22d1 U1845 ( .A1(n1072), .A2(\RegFilePlugin_regFile[13][16] ), .B1(n658), 
        .B2(\RegFilePlugin_regFile[10][16] ), .ZN(n1017) );
  aoi22d1 U1846 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][16] ), .B1(n1176), 
        .B2(\RegFilePlugin_regFile[2][16] ), .ZN(n1016) );
  aoi22d1 U1847 ( .A1(n1269), .A2(\RegFilePlugin_regFile[1][16] ), .B1(n1171), 
        .B2(\RegFilePlugin_regFile[11][16] ), .ZN(n1023) );
  aoi22d1 U1848 ( .A1(n988), .A2(\RegFilePlugin_regFile[28][16] ), .B1(n926), 
        .B2(\RegFilePlugin_regFile[0][16] ), .ZN(n1022) );
  aoi22d1 U1849 ( .A1(n867), .A2(\RegFilePlugin_regFile[24][16] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][16] ), .ZN(n1021) );
  aoi22d1 U1850 ( .A1(n1260), .A2(\RegFilePlugin_regFile[30][16] ), .B1(n1296), 
        .B2(\RegFilePlugin_regFile[12][16] ), .ZN(n1020) );
  aoi22d1 U1851 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][16] ), .B1(n1238), 
        .B2(\RegFilePlugin_regFile[4][16] ), .ZN(n1027) );
  aoi22d1 U1852 ( .A1(n1116), .A2(\RegFilePlugin_regFile[15][16] ), .B1(n1258), 
        .B2(\RegFilePlugin_regFile[21][16] ), .ZN(n1026) );
  aoi22d1 U1853 ( .A1(n1143), .A2(\RegFilePlugin_regFile[22][16] ), .B1(n1229), 
        .B2(\RegFilePlugin_regFile[9][16] ), .ZN(n1025) );
  aoi22d1 U1854 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][16] ), .B1(n757), 
        .B2(\RegFilePlugin_regFile[5][16] ), .ZN(n1024) );
  or04d0 U1855 ( .A1(n1031), .A2(n1030), .A3(n1029), .A4(n1028), .Z(N838) );
  aoi22d1 U1856 ( .A1(n1171), .A2(\RegFilePlugin_regFile[11][10] ), .B1(n1010), 
        .B2(\RegFilePlugin_regFile[16][10] ), .ZN(n1035) );
  aoi22d1 U1857 ( .A1(n1138), .A2(\RegFilePlugin_regFile[26][10] ), .B1(n1280), 
        .B2(\RegFilePlugin_regFile[3][10] ), .ZN(n1034) );
  aoi22d1 U1858 ( .A1(n1208), .A2(\RegFilePlugin_regFile[10][10] ), .B1(n988), 
        .B2(\RegFilePlugin_regFile[28][10] ), .ZN(n1033) );
  aoi22d1 U1859 ( .A1(n884), .A2(\RegFilePlugin_regFile[12][10] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][10] ), .ZN(n1032) );
  aoi22d1 U1860 ( .A1(n1275), .A2(\RegFilePlugin_regFile[6][10] ), .B1(n1270), 
        .B2(\RegFilePlugin_regFile[27][10] ), .ZN(n1039) );
  aoi22d1 U1861 ( .A1(n1253), .A2(\RegFilePlugin_regFile[7][10] ), .B1(n1271), 
        .B2(\RegFilePlugin_regFile[29][10] ), .ZN(n1038) );
  aoi22d1 U1862 ( .A1(n1072), .A2(\RegFilePlugin_regFile[13][10] ), .B1(n1166), 
        .B2(\RegFilePlugin_regFile[5][10] ), .ZN(n1037) );
  aoi22d1 U1863 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][10] ), .B1(n1148), 
        .B2(\RegFilePlugin_regFile[25][10] ), .ZN(n1036) );
  aoi22d1 U1864 ( .A1(n1143), .A2(\RegFilePlugin_regFile[22][10] ), .B1(n1209), 
        .B2(\RegFilePlugin_regFile[15][10] ), .ZN(n1043) );
  aoi22d1 U1865 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][10] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][10] ), .ZN(n1042) );
  aoi22d1 U1866 ( .A1(n1260), .A2(\RegFilePlugin_regFile[30][10] ), .B1(n841), 
        .B2(\RegFilePlugin_regFile[9][10] ), .ZN(n1041) );
  aoi22d1 U1867 ( .A1(n1259), .A2(\RegFilePlugin_regFile[1][10] ), .B1(n1238), 
        .B2(\RegFilePlugin_regFile[4][10] ), .ZN(n1040) );
  aoi22d1 U1868 ( .A1(n889), .A2(\RegFilePlugin_regFile[20][10] ), .B1(n1011), 
        .B2(\RegFilePlugin_regFile[31][10] ), .ZN(n1047) );
  aoi22d1 U1869 ( .A1(n1176), .A2(\RegFilePlugin_regFile[2][10] ), .B1(n1273), 
        .B2(\RegFilePlugin_regFile[24][10] ), .ZN(n1046) );
  aoi22d1 U1870 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][10] ), .B1(n1190), 
        .B2(\RegFilePlugin_regFile[19][10] ), .ZN(n1045) );
  aoi22d1 U1871 ( .A1(n1295), .A2(\RegFilePlugin_regFile[21][10] ), .B1(n779), 
        .B2(\RegFilePlugin_regFile[23][10] ), .ZN(n1044) );
  or04d0 U1872 ( .A1(n1051), .A2(n1050), .A3(n1049), .A4(n1048), .Z(N844) );
  aoi22d1 U1873 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][21] ), .B1(n779), 
        .B2(\RegFilePlugin_regFile[23][21] ), .ZN(n1055) );
  aoi22d1 U1874 ( .A1(n1116), .A2(\RegFilePlugin_regFile[15][21] ), .B1(n926), 
        .B2(\RegFilePlugin_regFile[0][21] ), .ZN(n1054) );
  aoi22d1 U1875 ( .A1(n1099), .A2(\RegFilePlugin_regFile[17][21] ), .B1(n842), 
        .B2(\RegFilePlugin_regFile[25][21] ), .ZN(n1053) );
  aoi22d1 U1876 ( .A1(n1275), .A2(\RegFilePlugin_regFile[6][21] ), .B1(n1252), 
        .B2(\RegFilePlugin_regFile[27][21] ), .ZN(n1052) );
  aoi22d1 U1877 ( .A1(n1222), .A2(\RegFilePlugin_regFile[20][21] ), .B1(n1297), 
        .B2(\RegFilePlugin_regFile[18][21] ), .ZN(n1059) );
  aoi22d1 U1878 ( .A1(n1072), .A2(\RegFilePlugin_regFile[13][21] ), .B1(n1176), 
        .B2(\RegFilePlugin_regFile[2][21] ), .ZN(n1058) );
  aoi22d1 U1879 ( .A1(n1138), .A2(\RegFilePlugin_regFile[26][21] ), .B1(n658), 
        .B2(\RegFilePlugin_regFile[10][21] ), .ZN(n1057) );
  aoi22d1 U1880 ( .A1(n884), .A2(\RegFilePlugin_regFile[12][21] ), .B1(n1011), 
        .B2(\RegFilePlugin_regFile[31][21] ), .ZN(n1056) );
  aoi22d1 U1881 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][21] ), .B1(n1273), 
        .B2(\RegFilePlugin_regFile[24][21] ), .ZN(n1063) );
  aoi22d1 U1882 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][21] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][21] ), .ZN(n1062) );
  aoi22d1 U1883 ( .A1(n1143), .A2(\RegFilePlugin_regFile[22][21] ), .B1(n1289), 
        .B2(\RegFilePlugin_regFile[7][21] ), .ZN(n1061) );
  aoi22d1 U1884 ( .A1(n1166), .A2(\RegFilePlugin_regFile[5][21] ), .B1(n1298), 
        .B2(\RegFilePlugin_regFile[28][21] ), .ZN(n1060) );
  aoi22d1 U1885 ( .A1(n1229), .A2(\RegFilePlugin_regFile[9][21] ), .B1(n1171), 
        .B2(\RegFilePlugin_regFile[11][21] ), .ZN(n1067) );
  aoi22d1 U1886 ( .A1(n1210), .A2(\RegFilePlugin_regFile[3][21] ), .B1(n1258), 
        .B2(\RegFilePlugin_regFile[21][21] ), .ZN(n1066) );
  aoi22d1 U1887 ( .A1(n1259), .A2(\RegFilePlugin_regFile[1][21] ), .B1(n1271), 
        .B2(\RegFilePlugin_regFile[29][21] ), .ZN(n1065) );
  aoi22d1 U1888 ( .A1(n1260), .A2(\RegFilePlugin_regFile[30][21] ), .B1(n1217), 
        .B2(\RegFilePlugin_regFile[4][21] ), .ZN(n1064) );
  or04d0 U1889 ( .A1(n1071), .A2(n1070), .A3(n1069), .A4(n1068), .Z(N833) );
  aoi22d1 U1890 ( .A1(n1138), .A2(\RegFilePlugin_regFile[26][4] ), .B1(n1222), 
        .B2(\RegFilePlugin_regFile[20][4] ), .ZN(n1077) );
  aoi22d1 U1891 ( .A1(n1072), .A2(\RegFilePlugin_regFile[13][4] ), .B1(n1238), 
        .B2(\RegFilePlugin_regFile[4][4] ), .ZN(n1076) );
  aoi22d1 U1892 ( .A1(n1073), .A2(\RegFilePlugin_regFile[2][4] ), .B1(n1208), 
        .B2(\RegFilePlugin_regFile[10][4] ), .ZN(n1075) );
  aoi22d1 U1893 ( .A1(n1253), .A2(\RegFilePlugin_regFile[7][4] ), .B1(n1171), 
        .B2(\RegFilePlugin_regFile[11][4] ), .ZN(n1074) );
  aoi22d1 U1894 ( .A1(n1099), .A2(\RegFilePlugin_regFile[17][4] ), .B1(n1209), 
        .B2(\RegFilePlugin_regFile[15][4] ), .ZN(n1081) );
  aoi22d1 U1895 ( .A1(n1294), .A2(\RegFilePlugin_regFile[8][4] ), .B1(n1143), 
        .B2(\RegFilePlugin_regFile[22][4] ), .ZN(n1080) );
  aoi22d1 U1896 ( .A1(n1270), .A2(\RegFilePlugin_regFile[27][4] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][4] ), .ZN(n1079) );
  aoi22d1 U1897 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][4] ), .B1(n1295), 
        .B2(\RegFilePlugin_regFile[21][4] ), .ZN(n1078) );
  aoi22d1 U1898 ( .A1(n653), .A2(\RegFilePlugin_regFile[30][4] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][4] ), .ZN(n1085) );
  aoi22d1 U1899 ( .A1(n1296), .A2(\RegFilePlugin_regFile[12][4] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][4] ), .ZN(n1084) );
  aoi22d1 U1900 ( .A1(n1273), .A2(\RegFilePlugin_regFile[24][4] ), .B1(n1281), 
        .B2(\RegFilePlugin_regFile[23][4] ), .ZN(n1083) );
  aoi22d1 U1901 ( .A1(n1269), .A2(\RegFilePlugin_regFile[1][4] ), .B1(n1166), 
        .B2(\RegFilePlugin_regFile[5][4] ), .ZN(n1082) );
  aoi22d1 U1902 ( .A1(n1275), .A2(\RegFilePlugin_regFile[6][4] ), .B1(n1011), 
        .B2(\RegFilePlugin_regFile[31][4] ), .ZN(n1089) );
  aoi22d1 U1903 ( .A1(n1271), .A2(\RegFilePlugin_regFile[29][4] ), .B1(n1229), 
        .B2(\RegFilePlugin_regFile[9][4] ), .ZN(n1088) );
  aoi22d1 U1904 ( .A1(n1148), .A2(\RegFilePlugin_regFile[25][4] ), .B1(n1280), 
        .B2(\RegFilePlugin_regFile[3][4] ), .ZN(n1087) );
  aoi22d1 U1905 ( .A1(n1190), .A2(\RegFilePlugin_regFile[19][4] ), .B1(n988), 
        .B2(\RegFilePlugin_regFile[28][4] ), .ZN(n1086) );
  or04d0 U1906 ( .A1(n1093), .A2(n1092), .A3(n1091), .A4(n1090), .Z(N850) );
  aoi22d1 U1907 ( .A1(n1094), .A2(\RegFilePlugin_regFile[29][12] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][12] ), .ZN(n1098) );
  aoi22d1 U1908 ( .A1(n842), .A2(\RegFilePlugin_regFile[25][12] ), .B1(n1273), 
        .B2(\RegFilePlugin_regFile[24][12] ), .ZN(n1097) );
  aoi22d1 U1909 ( .A1(n1253), .A2(\RegFilePlugin_regFile[7][12] ), .B1(n1166), 
        .B2(\RegFilePlugin_regFile[5][12] ), .ZN(n1096) );
  aoi22d1 U1910 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][12] ), .B1(n1208), 
        .B2(\RegFilePlugin_regFile[10][12] ), .ZN(n1095) );
  aoi22d1 U1911 ( .A1(n889), .A2(\RegFilePlugin_regFile[20][12] ), .B1(n1294), 
        .B2(\RegFilePlugin_regFile[8][12] ), .ZN(n1103) );
  aoi22d1 U1912 ( .A1(n1099), .A2(\RegFilePlugin_regFile[17][12] ), .B1(n1270), 
        .B2(\RegFilePlugin_regFile[27][12] ), .ZN(n1102) );
  aoi22d1 U1913 ( .A1(n1210), .A2(\RegFilePlugin_regFile[3][12] ), .B1(n779), 
        .B2(\RegFilePlugin_regFile[23][12] ), .ZN(n1101) );
  aoi22d1 U1914 ( .A1(n1297), .A2(\RegFilePlugin_regFile[18][12] ), .B1(n1229), 
        .B2(\RegFilePlugin_regFile[9][12] ), .ZN(n1100) );
  aoi22d1 U1915 ( .A1(n1288), .A2(\RegFilePlugin_regFile[22][12] ), .B1(n1295), 
        .B2(\RegFilePlugin_regFile[21][12] ), .ZN(n1107) );
  aoi22d1 U1916 ( .A1(n1072), .A2(\RegFilePlugin_regFile[13][12] ), .B1(n1238), 
        .B2(\RegFilePlugin_regFile[4][12] ), .ZN(n1106) );
  aoi22d1 U1917 ( .A1(n1190), .A2(\RegFilePlugin_regFile[19][12] ), .B1(n1250), 
        .B2(\RegFilePlugin_regFile[6][12] ), .ZN(n1105) );
  aoi22d1 U1918 ( .A1(n1116), .A2(\RegFilePlugin_regFile[15][12] ), .B1(n1272), 
        .B2(\RegFilePlugin_regFile[11][12] ), .ZN(n1104) );
  aoi22d1 U1919 ( .A1(n1073), .A2(\RegFilePlugin_regFile[2][12] ), .B1(n653), 
        .B2(\RegFilePlugin_regFile[30][12] ), .ZN(n1111) );
  aoi22d1 U1920 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][12] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][12] ), .ZN(n1110) );
  aoi22d1 U1921 ( .A1(n1259), .A2(\RegFilePlugin_regFile[1][12] ), .B1(n988), 
        .B2(\RegFilePlugin_regFile[28][12] ), .ZN(n1109) );
  aoi22d1 U1922 ( .A1(n884), .A2(\RegFilePlugin_regFile[12][12] ), .B1(n1010), 
        .B2(\RegFilePlugin_regFile[16][12] ), .ZN(n1108) );
  or04d0 U1923 ( .A1(n1115), .A2(n1114), .A3(n1113), .A4(n1112), .Z(N842) );
  aoi22d1 U1924 ( .A1(n1148), .A2(\RegFilePlugin_regFile[25][7] ), .B1(n1269), 
        .B2(\RegFilePlugin_regFile[1][7] ), .ZN(n1120) );
  aoi22d1 U1925 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][7] ), .B1(n1208), 
        .B2(\RegFilePlugin_regFile[10][7] ), .ZN(n1119) );
  aoi22d1 U1926 ( .A1(n1294), .A2(\RegFilePlugin_regFile[8][7] ), .B1(n1116), 
        .B2(\RegFilePlugin_regFile[15][7] ), .ZN(n1118) );
  aoi22d1 U1927 ( .A1(n1298), .A2(\RegFilePlugin_regFile[28][7] ), .B1(n1281), 
        .B2(\RegFilePlugin_regFile[23][7] ), .ZN(n1117) );
  aoi22d1 U1928 ( .A1(n867), .A2(\RegFilePlugin_regFile[24][7] ), .B1(n1010), 
        .B2(\RegFilePlugin_regFile[16][7] ), .ZN(n1125) );
  aoi22d1 U1929 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][7] ), .B1(n1275), 
        .B2(\RegFilePlugin_regFile[6][7] ), .ZN(n1124) );
  aoi22d1 U1930 ( .A1(n1244), .A2(\RegFilePlugin_regFile[13][7] ), .B1(n1166), 
        .B2(\RegFilePlugin_regFile[5][7] ), .ZN(n1123) );
  aoi22d1 U1931 ( .A1(n1288), .A2(\RegFilePlugin_regFile[22][7] ), .B1(n1271), 
        .B2(\RegFilePlugin_regFile[29][7] ), .ZN(n1122) );
  aoi22d1 U1932 ( .A1(n1280), .A2(\RegFilePlugin_regFile[3][7] ), .B1(n1272), 
        .B2(\RegFilePlugin_regFile[11][7] ), .ZN(n1129) );
  aoi22d1 U1933 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][7] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][7] ), .ZN(n1128) );
  aoi22d1 U1934 ( .A1(n1253), .A2(\RegFilePlugin_regFile[7][7] ), .B1(n1229), 
        .B2(\RegFilePlugin_regFile[9][7] ), .ZN(n1127) );
  aoi22d1 U1935 ( .A1(n1217), .A2(\RegFilePlugin_regFile[4][7] ), .B1(n884), 
        .B2(\RegFilePlugin_regFile[12][7] ), .ZN(n1126) );
  aoi22d1 U1936 ( .A1(n1176), .A2(\RegFilePlugin_regFile[2][7] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][7] ), .ZN(n1133) );
  aoi22d1 U1937 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][7] ), .B1(n653), 
        .B2(\RegFilePlugin_regFile[30][7] ), .ZN(n1132) );
  aoi22d1 U1938 ( .A1(n1222), .A2(\RegFilePlugin_regFile[20][7] ), .B1(n1295), 
        .B2(\RegFilePlugin_regFile[21][7] ), .ZN(n1131) );
  aoi22d1 U1939 ( .A1(n1252), .A2(\RegFilePlugin_regFile[27][7] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][7] ), .ZN(n1130) );
  or04d0 U1940 ( .A1(n1137), .A2(n1136), .A3(n1135), .A4(n1134), .Z(N847) );
  aoi22d1 U1941 ( .A1(n1072), .A2(\RegFilePlugin_regFile[13][8] ), .B1(n1250), 
        .B2(\RegFilePlugin_regFile[6][8] ), .ZN(n1142) );
  aoi22d1 U1942 ( .A1(n1138), .A2(\RegFilePlugin_regFile[26][8] ), .B1(n1297), 
        .B2(\RegFilePlugin_regFile[18][8] ), .ZN(n1141) );
  aoi22d1 U1943 ( .A1(n1260), .A2(\RegFilePlugin_regFile[30][8] ), .B1(n1217), 
        .B2(\RegFilePlugin_regFile[4][8] ), .ZN(n1140) );
  aoi22d1 U1944 ( .A1(n1298), .A2(\RegFilePlugin_regFile[28][8] ), .B1(n1010), 
        .B2(\RegFilePlugin_regFile[16][8] ), .ZN(n1139) );
  aoi22d1 U1945 ( .A1(n1190), .A2(\RegFilePlugin_regFile[19][8] ), .B1(n1222), 
        .B2(\RegFilePlugin_regFile[20][8] ), .ZN(n1147) );
  aoi22d1 U1946 ( .A1(n1143), .A2(\RegFilePlugin_regFile[22][8] ), .B1(n1253), 
        .B2(\RegFilePlugin_regFile[7][8] ), .ZN(n1146) );
  aoi22d1 U1947 ( .A1(n867), .A2(\RegFilePlugin_regFile[24][8] ), .B1(n1270), 
        .B2(\RegFilePlugin_regFile[27][8] ), .ZN(n1145) );
  aoi22d1 U1948 ( .A1(n658), .A2(\RegFilePlugin_regFile[10][8] ), .B1(n1272), 
        .B2(\RegFilePlugin_regFile[11][8] ), .ZN(n1144) );
  aoi22d1 U1949 ( .A1(n1148), .A2(\RegFilePlugin_regFile[25][8] ), .B1(n1271), 
        .B2(\RegFilePlugin_regFile[29][8] ), .ZN(n1152) );
  aoi22d1 U1950 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][8] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][8] ), .ZN(n1151) );
  aoi22d1 U1951 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][8] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][8] ), .ZN(n1150) );
  aoi22d1 U1952 ( .A1(n1099), .A2(\RegFilePlugin_regFile[17][8] ), .B1(n779), 
        .B2(\RegFilePlugin_regFile[23][8] ), .ZN(n1149) );
  aoi22d1 U1953 ( .A1(n1210), .A2(\RegFilePlugin_regFile[3][8] ), .B1(n1209), 
        .B2(\RegFilePlugin_regFile[15][8] ), .ZN(n1156) );
  aoi22d1 U1954 ( .A1(n1259), .A2(\RegFilePlugin_regFile[1][8] ), .B1(n1295), 
        .B2(\RegFilePlugin_regFile[21][8] ), .ZN(n1155) );
  aoi22d1 U1955 ( .A1(n1296), .A2(\RegFilePlugin_regFile[12][8] ), .B1(n841), 
        .B2(\RegFilePlugin_regFile[9][8] ), .ZN(n1154) );
  aoi22d1 U1956 ( .A1(n1073), .A2(\RegFilePlugin_regFile[2][8] ), .B1(n1166), 
        .B2(\RegFilePlugin_regFile[5][8] ), .ZN(n1153) );
  or04d0 U1957 ( .A1(n1160), .A2(n1159), .A3(n1158), .A4(n1157), .Z(N846) );
  aoi22d1 U1958 ( .A1(n1294), .A2(\RegFilePlugin_regFile[8][30] ), .B1(n1161), 
        .B2(\RegFilePlugin_regFile[6][30] ), .ZN(n1165) );
  aoi22d1 U1959 ( .A1(n1260), .A2(\RegFilePlugin_regFile[30][30] ), .B1(n1295), 
        .B2(\RegFilePlugin_regFile[21][30] ), .ZN(n1164) );
  aoi22d1 U1960 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][30] ), .B1(n842), 
        .B2(\RegFilePlugin_regFile[25][30] ), .ZN(n1163) );
  aoi22d1 U1961 ( .A1(n1244), .A2(\RegFilePlugin_regFile[13][30] ), .B1(n1010), 
        .B2(\RegFilePlugin_regFile[16][30] ), .ZN(n1162) );
  aoi22d1 U1962 ( .A1(n1208), .A2(\RegFilePlugin_regFile[10][30] ), .B1(n1166), 
        .B2(\RegFilePlugin_regFile[5][30] ), .ZN(n1170) );
  aoi22d1 U1963 ( .A1(n1222), .A2(\RegFilePlugin_regFile[20][30] ), .B1(n1259), 
        .B2(\RegFilePlugin_regFile[1][30] ), .ZN(n1169) );
  aoi22d1 U1964 ( .A1(n1252), .A2(\RegFilePlugin_regFile[27][30] ), .B1(n1281), 
        .B2(\RegFilePlugin_regFile[23][30] ), .ZN(n1168) );
  aoi22d1 U1965 ( .A1(n1238), .A2(\RegFilePlugin_regFile[4][30] ), .B1(n1297), 
        .B2(\RegFilePlugin_regFile[18][30] ), .ZN(n1167) );
  aoi22d1 U1966 ( .A1(n1282), .A2(\RegFilePlugin_regFile[14][30] ), .B1(n1171), 
        .B2(\RegFilePlugin_regFile[11][30] ), .ZN(n1175) );
  aoi22d1 U1967 ( .A1(n867), .A2(\RegFilePlugin_regFile[24][30] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][30] ), .ZN(n1174) );
  aoi22d1 U1968 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][30] ), .B1(n1280), 
        .B2(\RegFilePlugin_regFile[3][30] ), .ZN(n1173) );
  aoi22d1 U1969 ( .A1(n1271), .A2(\RegFilePlugin_regFile[29][30] ), .B1(n1209), 
        .B2(\RegFilePlugin_regFile[15][30] ), .ZN(n1172) );
  aoi22d1 U1970 ( .A1(n1288), .A2(\RegFilePlugin_regFile[22][30] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][30] ), .ZN(n1180) );
  aoi22d1 U1971 ( .A1(n1176), .A2(\RegFilePlugin_regFile[2][30] ), .B1(n988), 
        .B2(\RegFilePlugin_regFile[28][30] ), .ZN(n1179) );
  aoi22d1 U1972 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][30] ), .B1(n1296), 
        .B2(\RegFilePlugin_regFile[12][30] ), .ZN(n1178) );
  aoi22d1 U1973 ( .A1(n1289), .A2(\RegFilePlugin_regFile[7][30] ), .B1(n1229), 
        .B2(\RegFilePlugin_regFile[9][30] ), .ZN(n1177) );
  or04d0 U1974 ( .A1(n1184), .A2(n1183), .A3(n1182), .A4(n1181), .Z(N824) );
  aoi22d1 U1975 ( .A1(n1244), .A2(\RegFilePlugin_regFile[13][14] ), .B1(n1116), 
        .B2(\RegFilePlugin_regFile[15][14] ), .ZN(n1189) );
  aoi22d1 U1976 ( .A1(n1185), .A2(\RegFilePlugin_regFile[8][14] ), .B1(n1297), 
        .B2(\RegFilePlugin_regFile[18][14] ), .ZN(n1188) );
  aoi22d1 U1977 ( .A1(n1260), .A2(\RegFilePlugin_regFile[30][14] ), .B1(n1210), 
        .B2(\RegFilePlugin_regFile[3][14] ), .ZN(n1187) );
  aoi22d1 U1978 ( .A1(n1289), .A2(\RegFilePlugin_regFile[7][14] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][14] ), .ZN(n1186) );
  aoi22d1 U1979 ( .A1(n1099), .A2(\RegFilePlugin_regFile[17][14] ), .B1(n1190), 
        .B2(\RegFilePlugin_regFile[19][14] ), .ZN(n1194) );
  aoi22d1 U1980 ( .A1(n658), .A2(\RegFilePlugin_regFile[10][14] ), .B1(n884), 
        .B2(\RegFilePlugin_regFile[12][14] ), .ZN(n1193) );
  aoi22d1 U1981 ( .A1(n1270), .A2(\RegFilePlugin_regFile[27][14] ), .B1(n841), 
        .B2(\RegFilePlugin_regFile[9][14] ), .ZN(n1192) );
  aoi22d1 U1982 ( .A1(n1250), .A2(\RegFilePlugin_regFile[6][14] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][14] ), .ZN(n1191) );
  aoi22d1 U1983 ( .A1(n779), .A2(\RegFilePlugin_regFile[23][14] ), .B1(n1011), 
        .B2(\RegFilePlugin_regFile[31][14] ), .ZN(n1199) );
  aoi22d1 U1984 ( .A1(n1288), .A2(\RegFilePlugin_regFile[22][14] ), .B1(n1273), 
        .B2(\RegFilePlugin_regFile[24][14] ), .ZN(n1198) );
  aoi22d1 U1985 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][14] ), .B1(n757), 
        .B2(\RegFilePlugin_regFile[5][14] ), .ZN(n1197) );
  aoi22d1 U1986 ( .A1(n1258), .A2(\RegFilePlugin_regFile[21][14] ), .B1(n1272), 
        .B2(\RegFilePlugin_regFile[11][14] ), .ZN(n1196) );
  aoi22d1 U1987 ( .A1(n1222), .A2(\RegFilePlugin_regFile[20][14] ), .B1(n1282), 
        .B2(\RegFilePlugin_regFile[14][14] ), .ZN(n1203) );
  aoi22d1 U1988 ( .A1(n1217), .A2(\RegFilePlugin_regFile[4][14] ), .B1(n1271), 
        .B2(\RegFilePlugin_regFile[29][14] ), .ZN(n1202) );
  aoi22d1 U1989 ( .A1(n842), .A2(\RegFilePlugin_regFile[25][14] ), .B1(n1298), 
        .B2(\RegFilePlugin_regFile[28][14] ), .ZN(n1201) );
  aoi22d1 U1990 ( .A1(n1073), .A2(\RegFilePlugin_regFile[2][14] ), .B1(n1269), 
        .B2(\RegFilePlugin_regFile[1][14] ), .ZN(n1200) );
  or04d0 U1991 ( .A1(n1207), .A2(n1206), .A3(n1205), .A4(n1204), .Z(N840) );
  aoi22d1 U1992 ( .A1(n1288), .A2(\RegFilePlugin_regFile[22][23] ), .B1(n1208), 
        .B2(\RegFilePlugin_regFile[10][23] ), .ZN(n1214) );
  aoi22d1 U1993 ( .A1(n1195), .A2(\RegFilePlugin_regFile[26][23] ), .B1(n842), 
        .B2(\RegFilePlugin_regFile[25][23] ), .ZN(n1213) );
  aoi22d1 U1994 ( .A1(n1210), .A2(\RegFilePlugin_regFile[3][23] ), .B1(n1209), 
        .B2(\RegFilePlugin_regFile[15][23] ), .ZN(n1212) );
  aoi22d1 U1995 ( .A1(n1176), .A2(\RegFilePlugin_regFile[2][23] ), .B1(n1252), 
        .B2(\RegFilePlugin_regFile[27][23] ), .ZN(n1211) );
  aoi22d1 U1996 ( .A1(n1296), .A2(\RegFilePlugin_regFile[12][23] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][23] ), .ZN(n1221) );
  aoi22d1 U1997 ( .A1(n1216), .A2(\RegFilePlugin_regFile[7][23] ), .B1(n1275), 
        .B2(\RegFilePlugin_regFile[6][23] ), .ZN(n1220) );
  aoi22d1 U1998 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][23] ), .B1(n1217), 
        .B2(\RegFilePlugin_regFile[4][23] ), .ZN(n1219) );
  aoi22d1 U1999 ( .A1(n1072), .A2(\RegFilePlugin_regFile[13][23] ), .B1(n1298), 
        .B2(\RegFilePlugin_regFile[28][23] ), .ZN(n1218) );
  aoi22d1 U2000 ( .A1(n1222), .A2(\RegFilePlugin_regFile[20][23] ), .B1(n1281), 
        .B2(\RegFilePlugin_regFile[23][23] ), .ZN(n1227) );
  aoi22d1 U2001 ( .A1(n1099), .A2(\RegFilePlugin_regFile[17][23] ), .B1(n1094), 
        .B2(\RegFilePlugin_regFile[29][23] ), .ZN(n1226) );
  aoi22d1 U2002 ( .A1(n1273), .A2(\RegFilePlugin_regFile[24][23] ), .B1(n1223), 
        .B2(\RegFilePlugin_regFile[18][23] ), .ZN(n1225) );
  aoi22d1 U2003 ( .A1(n1282), .A2(\RegFilePlugin_regFile[14][23] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][23] ), .ZN(n1224) );
  aoi22d1 U2004 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][23] ), .B1(n1258), 
        .B2(\RegFilePlugin_regFile[21][23] ), .ZN(n1233) );
  aoi22d1 U2005 ( .A1(n653), .A2(\RegFilePlugin_regFile[30][23] ), .B1(n757), 
        .B2(\RegFilePlugin_regFile[5][23] ), .ZN(n1232) );
  aoi22d1 U2006 ( .A1(n1269), .A2(\RegFilePlugin_regFile[1][23] ), .B1(n1272), 
        .B2(\RegFilePlugin_regFile[11][23] ), .ZN(n1231) );
  aoi22d1 U2007 ( .A1(n1229), .A2(\RegFilePlugin_regFile[9][23] ), .B1(n1228), 
        .B2(\RegFilePlugin_regFile[31][23] ), .ZN(n1230) );
  or04d0 U2008 ( .A1(n1237), .A2(n1236), .A3(n1235), .A4(n1234), .Z(N831) );
  aoi22d1 U2009 ( .A1(n1272), .A2(\RegFilePlugin_regFile[11][15] ), .B1(n1281), 
        .B2(\RegFilePlugin_regFile[23][15] ), .ZN(n1243) );
  aoi22d1 U2010 ( .A1(n1238), .A2(\RegFilePlugin_regFile[4][15] ), .B1(n867), 
        .B2(\RegFilePlugin_regFile[24][15] ), .ZN(n1242) );
  aoi22d1 U2011 ( .A1(n1239), .A2(\RegFilePlugin_regFile[8][15] ), .B1(n1271), 
        .B2(\RegFilePlugin_regFile[29][15] ), .ZN(n1241) );
  aoi22d1 U2012 ( .A1(n1138), .A2(\RegFilePlugin_regFile[26][15] ), .B1(n1116), 
        .B2(\RegFilePlugin_regFile[15][15] ), .ZN(n1240) );
  aoi22d1 U2013 ( .A1(n1244), .A2(\RegFilePlugin_regFile[13][15] ), .B1(n1296), 
        .B2(\RegFilePlugin_regFile[12][15] ), .ZN(n1249) );
  aoi22d1 U2014 ( .A1(n1245), .A2(\RegFilePlugin_regFile[14][15] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][15] ), .ZN(n1248) );
  aoi22d1 U2015 ( .A1(n1297), .A2(\RegFilePlugin_regFile[18][15] ), .B1(n1011), 
        .B2(\RegFilePlugin_regFile[31][15] ), .ZN(n1247) );
  aoi22d1 U2016 ( .A1(n1143), .A2(\RegFilePlugin_regFile[22][15] ), .B1(n1298), 
        .B2(\RegFilePlugin_regFile[28][15] ), .ZN(n1246) );
  aoi22d1 U2017 ( .A1(n1176), .A2(\RegFilePlugin_regFile[2][15] ), .B1(n1250), 
        .B2(\RegFilePlugin_regFile[6][15] ), .ZN(n1257) );
  aoi22d1 U2018 ( .A1(n1251), .A2(\RegFilePlugin_regFile[17][15] ), .B1(n1210), 
        .B2(\RegFilePlugin_regFile[3][15] ), .ZN(n1256) );
  aoi22d1 U2019 ( .A1(n889), .A2(\RegFilePlugin_regFile[20][15] ), .B1(n1252), 
        .B2(\RegFilePlugin_regFile[27][15] ), .ZN(n1255) );
  aoi22d1 U2020 ( .A1(n1253), .A2(\RegFilePlugin_regFile[7][15] ), .B1(n757), 
        .B2(\RegFilePlugin_regFile[5][15] ), .ZN(n1254) );
  aoi22d1 U2021 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][15] ), .B1(n1229), 
        .B2(\RegFilePlugin_regFile[9][15] ), .ZN(n1264) );
  aoi22d1 U2022 ( .A1(n1259), .A2(\RegFilePlugin_regFile[1][15] ), .B1(n1258), 
        .B2(\RegFilePlugin_regFile[21][15] ), .ZN(n1263) );
  aoi22d1 U2023 ( .A1(n842), .A2(\RegFilePlugin_regFile[25][15] ), .B1(n1208), 
        .B2(\RegFilePlugin_regFile[10][15] ), .ZN(n1262) );
  aoi22d1 U2024 ( .A1(n1260), .A2(\RegFilePlugin_regFile[30][15] ), .B1(n1215), 
        .B2(\RegFilePlugin_regFile[0][15] ), .ZN(n1261) );
  or04d0 U2025 ( .A1(n1268), .A2(n1267), .A3(n1266), .A4(n1265), .Z(N839) );
  aoi22d1 U2026 ( .A1(n1269), .A2(\RegFilePlugin_regFile[1][18] ), .B1(n1238), 
        .B2(\RegFilePlugin_regFile[4][18] ), .ZN(n1279) );
  aoi22d1 U2027 ( .A1(n1271), .A2(\RegFilePlugin_regFile[29][18] ), .B1(n1270), 
        .B2(\RegFilePlugin_regFile[27][18] ), .ZN(n1278) );
  aoi22d1 U2028 ( .A1(n1273), .A2(\RegFilePlugin_regFile[24][18] ), .B1(n1272), 
        .B2(\RegFilePlugin_regFile[11][18] ), .ZN(n1277) );
  aoi22d1 U2029 ( .A1(n1275), .A2(\RegFilePlugin_regFile[6][18] ), .B1(n1274), 
        .B2(\RegFilePlugin_regFile[16][18] ), .ZN(n1276) );
  aoi22d1 U2030 ( .A1(n889), .A2(\RegFilePlugin_regFile[20][18] ), .B1(n1280), 
        .B2(\RegFilePlugin_regFile[3][18] ), .ZN(n1286) );
  aoi22d1 U2031 ( .A1(n1138), .A2(\RegFilePlugin_regFile[26][18] ), .B1(n757), 
        .B2(\RegFilePlugin_regFile[5][18] ), .ZN(n1285) );
  aoi22d1 U2032 ( .A1(n1282), .A2(\RegFilePlugin_regFile[14][18] ), .B1(n1281), 
        .B2(\RegFilePlugin_regFile[23][18] ), .ZN(n1284) );
  aoi22d1 U2033 ( .A1(n1072), .A2(\RegFilePlugin_regFile[13][18] ), .B1(n841), 
        .B2(\RegFilePlugin_regFile[9][18] ), .ZN(n1283) );
  aoi22d1 U2034 ( .A1(n1287), .A2(\RegFilePlugin_regFile[19][18] ), .B1(n842), 
        .B2(\RegFilePlugin_regFile[25][18] ), .ZN(n1293) );
  aoi22d1 U2035 ( .A1(n1073), .A2(\RegFilePlugin_regFile[2][18] ), .B1(n1288), 
        .B2(\RegFilePlugin_regFile[22][18] ), .ZN(n1292) );
  aoi22d1 U2036 ( .A1(n658), .A2(\RegFilePlugin_regFile[10][18] ), .B1(n653), 
        .B2(\RegFilePlugin_regFile[30][18] ), .ZN(n1291) );
  aoi22d1 U2037 ( .A1(n1289), .A2(\RegFilePlugin_regFile[7][18] ), .B1(n1116), 
        .B2(\RegFilePlugin_regFile[15][18] ), .ZN(n1290) );
  aoi22d1 U2038 ( .A1(n1294), .A2(\RegFilePlugin_regFile[8][18] ), .B1(n1011), 
        .B2(\RegFilePlugin_regFile[31][18] ), .ZN(n1302) );
  aoi22d1 U2039 ( .A1(n1295), .A2(\RegFilePlugin_regFile[21][18] ), .B1(n926), 
        .B2(\RegFilePlugin_regFile[0][18] ), .ZN(n1301) );
  aoi22d1 U2040 ( .A1(n1297), .A2(\RegFilePlugin_regFile[18][18] ), .B1(n1296), 
        .B2(\RegFilePlugin_regFile[12][18] ), .ZN(n1300) );
  aoi22d1 U2041 ( .A1(n1099), .A2(\RegFilePlugin_regFile[17][18] ), .B1(n1298), 
        .B2(\RegFilePlugin_regFile[28][18] ), .ZN(n1299) );
  or04d0 U2042 ( .A1(n1306), .A2(n1305), .A3(n1304), .A4(n1303), .Z(N836) );
  aoi22d1 U2043 ( .A1(n3818), .A2(IBusCachedPlugin_cache_io_cpu_fetch_data[20]), .B1(\_zz__zz_decode_ENV_CTRL_2_1[20] ), .B2(n2374), .ZN(n1308) );
  inv0d0 U2044 ( .I(IBusCachedPlugin_cache_io_cpu_fetch_data[21]), .ZN(n6562)
         );
  aoi22d1 U2045 ( .A1(n3818), .A2(n6562), .B1(n2616), .B2(n2374), .ZN(n1309)
         );
  aoi22d1 U2046 ( .A1(n3818), .A2(IBusCachedPlugin_cache_io_cpu_fetch_data[23]), .B1(decode_INSTRUCTION_23), .B2(n2374), .ZN(n1316) );
  inv0d0 U2047 ( .I(IBusCachedPlugin_cache_io_cpu_fetch_data[24]), .ZN(n6523)
         );
  aoi22d1 U2048 ( .A1(n3818), .A2(n6523), .B1(n2613), .B2(n2374), .ZN(n1313)
         );
  aoi22d1 U2049 ( .A1(n3818), .A2(IBusCachedPlugin_cache_io_cpu_fetch_data[22]), .B1(decode_INSTRUCTION_22), .B2(n2374), .ZN(n1314) );
  inv0d0 U2050 ( .I(n1314), .ZN(n1307) );
  nr02d1 U2051 ( .A1(n1340), .A2(n1325), .ZN(n1628) );
  buffd1 U2052 ( .I(n1628), .Z(n2032) );
  inv0d0 U2053 ( .I(n1309), .ZN(n1311) );
  inv0d0 U2054 ( .I(n1313), .ZN(n1312) );
  inv0d0 U2055 ( .I(n1316), .ZN(n1323) );
  nr02d1 U2056 ( .A1(n1331), .A2(n1336), .ZN(n1735) );
  buffd1 U2057 ( .I(n1735), .Z(n2020) );
  aoi22d1 U2058 ( .A1(\RegFilePlugin_regFile[2][28] ), .A2(n2032), .B1(
        \RegFilePlugin_regFile[24][28] ), .B2(n2020), .ZN(n1320) );
  inv0d0 U2059 ( .I(n1308), .ZN(n1310) );
  nr02d1 U2060 ( .A1(n1341), .A2(n1325), .ZN(n1816) );
  nr02d1 U2061 ( .A1(n1344), .A2(n1339), .ZN(n1377) );
  buffd1 U2062 ( .I(n1377), .Z(n1931) );
  aoi22d1 U2063 ( .A1(\RegFilePlugin_regFile[3][28] ), .A2(n1816), .B1(
        \RegFilePlugin_regFile[21][28] ), .B2(n1931), .ZN(n1319) );
  nr02d1 U2064 ( .A1(n1331), .A2(n1339), .ZN(n1387) );
  buffd1 U2065 ( .I(n1387), .Z(n2006) );
  nr02d0 U2066 ( .A1(n1314), .A2(n1313), .ZN(n1324) );
  nr02d1 U2067 ( .A1(n1337), .A2(n1341), .ZN(n1543) );
  buffd1 U2068 ( .I(n1543), .Z(n1925) );
  aoi22d1 U2069 ( .A1(\RegFilePlugin_regFile[20][28] ), .A2(n2006), .B1(
        \RegFilePlugin_regFile[7][28] ), .B2(n1925), .ZN(n1318) );
  nr02d1 U2070 ( .A1(n1331), .A2(n1342), .ZN(n1671) );
  buffd1 U2071 ( .I(n1671), .Z(n1975) );
  nr02d1 U2072 ( .A1(n1331), .A2(n1337), .ZN(n1879) );
  buffd1 U2073 ( .I(n1879), .Z(n2004) );
  aoi22d1 U2074 ( .A1(\RegFilePlugin_regFile[16][28] ), .A2(n1975), .B1(
        \RegFilePlugin_regFile[4][28] ), .B2(n2004), .ZN(n1317) );
  nr02d1 U2075 ( .A1(n1336), .A2(n1340), .ZN(n1649) );
  buffd1 U2076 ( .I(n1649), .Z(n2015) );
  nr02d1 U2077 ( .A1(n1343), .A2(n1341), .ZN(n1901) );
  buffd1 U2078 ( .I(n1901), .Z(n2013) );
  aoi22d1 U2079 ( .A1(\RegFilePlugin_regFile[26][28] ), .A2(n2015), .B1(
        \RegFilePlugin_regFile[11][28] ), .B2(n2013), .ZN(n1329) );
  nr02d1 U2080 ( .A1(n1339), .A2(n1341), .ZN(n1544) );
  buffd1 U2081 ( .I(n1544), .Z(n2021) );
  nr02d1 U2082 ( .A1(n1344), .A2(n1325), .ZN(n1692) );
  buffd1 U2083 ( .I(n1692), .Z(n2012) );
  aoi22d1 U2084 ( .A1(\RegFilePlugin_regFile[23][28] ), .A2(n2021), .B1(
        \RegFilePlugin_regFile[1][28] ), .B2(n2012), .ZN(n1328) );
  nr02d1 U2085 ( .A1(n1330), .A2(n1344), .ZN(n1501) );
  buffd1 U2086 ( .I(n1501), .Z(n1974) );
  buffd1 U2087 ( .I(n1378), .Z(n1916) );
  aoi22d1 U2088 ( .A1(\RegFilePlugin_regFile[29][28] ), .A2(n1974), .B1(
        \RegFilePlugin_regFile[14][28] ), .B2(n1916), .ZN(n1327) );
  nr02d1 U2089 ( .A1(n1331), .A2(n1325), .ZN(n1585) );
  buffd1 U2090 ( .I(n1585), .Z(n2030) );
  buffd1 U2091 ( .I(n1697), .Z(n2023) );
  aoi22d1 U2092 ( .A1(\RegFilePlugin_regFile[0][28] ), .A2(n2030), .B1(
        \RegFilePlugin_regFile[15][28] ), .B2(n2023), .ZN(n1326) );
  nr02d1 U2093 ( .A1(n1330), .A2(n1341), .ZN(n1417) );
  buffd1 U2094 ( .I(n1417), .Z(n1942) );
  nr02d1 U2095 ( .A1(n1340), .A2(n1330), .ZN(n1837) );
  buffd1 U2096 ( .I(n1837), .Z(n1987) );
  aoi22d1 U2097 ( .A1(\RegFilePlugin_regFile[31][28] ), .A2(n1942), .B1(
        \RegFilePlugin_regFile[30][28] ), .B2(n1987), .ZN(n1335) );
  nr02d1 U2098 ( .A1(n1340), .A2(n1343), .ZN(n1416) );
  buffd1 U2099 ( .I(n1416), .Z(n1993) );
  nr02d1 U2100 ( .A1(n1331), .A2(n1343), .ZN(n1670) );
  buffd1 U2101 ( .I(n1670), .Z(n1902) );
  aoi22d1 U2102 ( .A1(\RegFilePlugin_regFile[10][28] ), .A2(n1993), .B1(
        \RegFilePlugin_regFile[8][28] ), .B2(n1902), .ZN(n1334) );
  nr02d1 U2103 ( .A1(n1340), .A2(n1342), .ZN(n1952) );
  buffd1 U2104 ( .I(n1952), .Z(n1937) );
  buffd1 U2105 ( .I(n2005), .Z(n1953) );
  aoi22d1 U2106 ( .A1(\RegFilePlugin_regFile[18][28] ), .A2(n1937), .B1(
        \RegFilePlugin_regFile[17][28] ), .B2(n1953), .ZN(n1333) );
  buffd1 U2107 ( .I(n1463), .Z(n2031) );
  nr02d1 U2108 ( .A1(n1331), .A2(n1330), .ZN(n1903) );
  buffd1 U2109 ( .I(n1903), .Z(n1892) );
  aoi22d1 U2110 ( .A1(\RegFilePlugin_regFile[12][28] ), .A2(n2031), .B1(
        \RegFilePlugin_regFile[28][28] ), .B2(n1892), .ZN(n1332) );
  nr02d1 U2111 ( .A1(n1337), .A2(n1344), .ZN(n1606) );
  buffd1 U2112 ( .I(n1606), .Z(n1982) );
  nr02d1 U2113 ( .A1(n1336), .A2(n1341), .ZN(n1718) );
  buffd1 U2114 ( .I(n1718), .Z(n2033) );
  aoi22d1 U2115 ( .A1(\RegFilePlugin_regFile[5][28] ), .A2(n1982), .B1(
        \RegFilePlugin_regFile[27][28] ), .B2(n2033), .ZN(n1348) );
  nr02d1 U2116 ( .A1(n1336), .A2(n1344), .ZN(n1607) );
  buffd1 U2117 ( .I(n1607), .Z(n1926) );
  nr02d1 U2118 ( .A1(n1337), .A2(n1340), .ZN(n1522) );
  buffd1 U2119 ( .I(n1522), .Z(n1943) );
  aoi22d1 U2120 ( .A1(\RegFilePlugin_regFile[25][28] ), .A2(n1926), .B1(
        \RegFilePlugin_regFile[6][28] ), .B2(n1943), .ZN(n1347) );
  nr02d1 U2121 ( .A1(n1344), .A2(n1338), .ZN(n1932) );
  buffd1 U2122 ( .I(n1932), .Z(n2025) );
  buffd1 U2123 ( .I(n1472), .Z(n2014) );
  aoi22d1 U2124 ( .A1(\RegFilePlugin_regFile[13][28] ), .A2(n2025), .B1(
        \RegFilePlugin_regFile[22][28] ), .B2(n2014), .ZN(n1346) );
  nr02d1 U2125 ( .A1(n1342), .A2(n1341), .ZN(n1458) );
  buffd1 U2126 ( .I(n1458), .Z(n2024) );
  nr02d1 U2127 ( .A1(n1344), .A2(n1343), .ZN(n1858) );
  buffd1 U2128 ( .I(n1858), .Z(n2011) );
  aoi22d1 U2129 ( .A1(\RegFilePlugin_regFile[19][28] ), .A2(n2024), .B1(
        \RegFilePlugin_regFile[9][28] ), .B2(n2011), .ZN(n1345) );
  or04d0 U2130 ( .A1(n1352), .A2(n1351), .A3(n1350), .A4(n1349), .Z(N859) );
  buffd1 U2131 ( .I(n1816), .Z(n2022) );
  aoi22d1 U2132 ( .A1(\RegFilePlugin_regFile[1][9] ), .A2(n2012), .B1(
        \RegFilePlugin_regFile[3][9] ), .B2(n2022), .ZN(n1356) );
  aoi22d1 U2133 ( .A1(\RegFilePlugin_regFile[6][9] ), .A2(n1522), .B1(
        \RegFilePlugin_regFile[27][9] ), .B2(n1718), .ZN(n1355) );
  buffd1 U2134 ( .I(n1378), .Z(n2003) );
  aoi22d1 U2135 ( .A1(\RegFilePlugin_regFile[14][9] ), .A2(n2003), .B1(
        \RegFilePlugin_regFile[9][9] ), .B2(n2011), .ZN(n1354) );
  aoi22d1 U2136 ( .A1(\RegFilePlugin_regFile[10][9] ), .A2(n1993), .B1(
        \RegFilePlugin_regFile[24][9] ), .B2(n2020), .ZN(n1353) );
  aoi22d1 U2137 ( .A1(\RegFilePlugin_regFile[16][9] ), .A2(n1975), .B1(
        \RegFilePlugin_regFile[29][9] ), .B2(n1501), .ZN(n1360) );
  buffd1 U2138 ( .I(n2005), .Z(n1976) );
  aoi22d1 U2139 ( .A1(\RegFilePlugin_regFile[20][9] ), .A2(n1387), .B1(
        \RegFilePlugin_regFile[17][9] ), .B2(n1976), .ZN(n1359) );
  aoi22d1 U2140 ( .A1(\RegFilePlugin_regFile[4][9] ), .A2(n1879), .B1(
        \RegFilePlugin_regFile[18][9] ), .B2(n1952), .ZN(n1358) );
  aoi22d1 U2141 ( .A1(\RegFilePlugin_regFile[28][9] ), .A2(n1903), .B1(
        \RegFilePlugin_regFile[19][9] ), .B2(n1458), .ZN(n1357) );
  buffd1 U2142 ( .I(n1697), .Z(n1994) );
  aoi22d1 U2143 ( .A1(\RegFilePlugin_regFile[26][9] ), .A2(n1649), .B1(
        \RegFilePlugin_regFile[15][9] ), .B2(n1994), .ZN(n1364) );
  aoi22d1 U2144 ( .A1(\RegFilePlugin_regFile[8][9] ), .A2(n1670), .B1(
        \RegFilePlugin_regFile[22][9] ), .B2(n2014), .ZN(n1363) );
  aoi22d1 U2145 ( .A1(\RegFilePlugin_regFile[11][9] ), .A2(n1901), .B1(
        \RegFilePlugin_regFile[0][9] ), .B2(n1585), .ZN(n1362) );
  aoi22d1 U2146 ( .A1(\RegFilePlugin_regFile[30][9] ), .A2(n1987), .B1(
        \RegFilePlugin_regFile[31][9] ), .B2(n1942), .ZN(n1361) );
  aoi22d1 U2147 ( .A1(\RegFilePlugin_regFile[12][9] ), .A2(n2031), .B1(
        \RegFilePlugin_regFile[21][9] ), .B2(n1931), .ZN(n1368) );
  aoi22d1 U2148 ( .A1(\RegFilePlugin_regFile[5][9] ), .A2(n1982), .B1(
        \RegFilePlugin_regFile[2][9] ), .B2(n1628), .ZN(n1367) );
  aoi22d1 U2149 ( .A1(\RegFilePlugin_regFile[23][9] ), .A2(n2021), .B1(
        \RegFilePlugin_regFile[7][9] ), .B2(n1925), .ZN(n1366) );
  aoi22d1 U2150 ( .A1(\RegFilePlugin_regFile[25][9] ), .A2(n1607), .B1(
        \RegFilePlugin_regFile[13][9] ), .B2(n2025), .ZN(n1365) );
  or04d0 U2151 ( .A1(n1372), .A2(n1371), .A3(n1370), .A4(n1369), .Z(N878) );
  aoi22d1 U2152 ( .A1(\RegFilePlugin_regFile[28][0] ), .A2(n1903), .B1(
        \RegFilePlugin_regFile[11][0] ), .B2(n1901), .ZN(n1376) );
  aoi22d1 U2153 ( .A1(\RegFilePlugin_regFile[23][0] ), .A2(n1544), .B1(
        \RegFilePlugin_regFile[31][0] ), .B2(n1417), .ZN(n1375) );
  aoi22d1 U2154 ( .A1(\RegFilePlugin_regFile[5][0] ), .A2(n1606), .B1(
        \RegFilePlugin_regFile[25][0] ), .B2(n1607), .ZN(n1374) );
  aoi22d1 U2155 ( .A1(\RegFilePlugin_regFile[9][0] ), .A2(n1858), .B1(
        \RegFilePlugin_regFile[30][0] ), .B2(n1987), .ZN(n1373) );
  aoi22d1 U2156 ( .A1(\RegFilePlugin_regFile[21][0] ), .A2(n1377), .B1(
        \RegFilePlugin_regFile[10][0] ), .B2(n1993), .ZN(n1382) );
  aoi22d1 U2157 ( .A1(\RegFilePlugin_regFile[8][0] ), .A2(n1902), .B1(
        \RegFilePlugin_regFile[26][0] ), .B2(n2015), .ZN(n1381) );
  aoi22d1 U2158 ( .A1(\RegFilePlugin_regFile[0][0] ), .A2(n1585), .B1(
        \RegFilePlugin_regFile[14][0] ), .B2(n1378), .ZN(n1380) );
  aoi22d1 U2159 ( .A1(\RegFilePlugin_regFile[27][0] ), .A2(n1718), .B1(
        \RegFilePlugin_regFile[1][0] ), .B2(n2012), .ZN(n1379) );
  aoi22d1 U2160 ( .A1(\RegFilePlugin_regFile[22][0] ), .A2(n2014), .B1(
        \RegFilePlugin_regFile[18][0] ), .B2(n1937), .ZN(n1386) );
  aoi22d1 U2161 ( .A1(\RegFilePlugin_regFile[16][0] ), .A2(n1975), .B1(
        \RegFilePlugin_regFile[7][0] ), .B2(n1543), .ZN(n1385) );
  aoi22d1 U2162 ( .A1(\RegFilePlugin_regFile[29][0] ), .A2(n1974), .B1(
        \RegFilePlugin_regFile[15][0] ), .B2(n1994), .ZN(n1384) );
  aoi22d1 U2163 ( .A1(\RegFilePlugin_regFile[6][0] ), .A2(n1522), .B1(
        \RegFilePlugin_regFile[3][0] ), .B2(n2022), .ZN(n1383) );
  aoi22d1 U2164 ( .A1(\RegFilePlugin_regFile[12][0] ), .A2(n2031), .B1(
        \RegFilePlugin_regFile[17][0] ), .B2(n1953), .ZN(n1391) );
  aoi22d1 U2165 ( .A1(\RegFilePlugin_regFile[24][0] ), .A2(n1735), .B1(
        \RegFilePlugin_regFile[2][0] ), .B2(n1628), .ZN(n1390) );
  aoi22d1 U2166 ( .A1(\RegFilePlugin_regFile[13][0] ), .A2(n1932), .B1(
        \RegFilePlugin_regFile[4][0] ), .B2(n2004), .ZN(n1389) );
  aoi22d1 U2167 ( .A1(\RegFilePlugin_regFile[20][0] ), .A2(n1387), .B1(
        \RegFilePlugin_regFile[19][0] ), .B2(n2024), .ZN(n1388) );
  or04d0 U2168 ( .A1(n1395), .A2(n1394), .A3(n1393), .A4(n1392), .Z(N887) );
  aoi22d1 U2169 ( .A1(\RegFilePlugin_regFile[4][27] ), .A2(n1879), .B1(
        \RegFilePlugin_regFile[12][27] ), .B2(n2031), .ZN(n1399) );
  aoi22d1 U2170 ( .A1(\RegFilePlugin_regFile[1][27] ), .A2(n1692), .B1(
        \RegFilePlugin_regFile[3][27] ), .B2(n1816), .ZN(n1398) );
  aoi22d1 U2171 ( .A1(\RegFilePlugin_regFile[30][27] ), .A2(n1987), .B1(
        \RegFilePlugin_regFile[27][27] ), .B2(n2033), .ZN(n1397) );
  aoi22d1 U2172 ( .A1(\RegFilePlugin_regFile[24][27] ), .A2(n2020), .B1(
        \RegFilePlugin_regFile[7][27] ), .B2(n1925), .ZN(n1396) );
  aoi22d1 U2173 ( .A1(\RegFilePlugin_regFile[20][27] ), .A2(n2006), .B1(
        \RegFilePlugin_regFile[14][27] ), .B2(n1916), .ZN(n1403) );
  aoi22d1 U2174 ( .A1(\RegFilePlugin_regFile[6][27] ), .A2(n1943), .B1(
        \RegFilePlugin_regFile[9][27] ), .B2(n2011), .ZN(n1402) );
  aoi22d1 U2175 ( .A1(\RegFilePlugin_regFile[5][27] ), .A2(n1606), .B1(
        \RegFilePlugin_regFile[22][27] ), .B2(n2014), .ZN(n1401) );
  aoi22d1 U2176 ( .A1(\RegFilePlugin_regFile[11][27] ), .A2(n1901), .B1(
        \RegFilePlugin_regFile[19][27] ), .B2(n1458), .ZN(n1400) );
  aoi22d1 U2177 ( .A1(\RegFilePlugin_regFile[28][27] ), .A2(n1903), .B1(
        \RegFilePlugin_regFile[18][27] ), .B2(n1952), .ZN(n1407) );
  aoi22d1 U2178 ( .A1(\RegFilePlugin_regFile[13][27] ), .A2(n2025), .B1(
        \RegFilePlugin_regFile[21][27] ), .B2(n1931), .ZN(n1406) );
  aoi22d1 U2179 ( .A1(\RegFilePlugin_regFile[25][27] ), .A2(n1926), .B1(
        \RegFilePlugin_regFile[31][27] ), .B2(n1942), .ZN(n1405) );
  aoi22d1 U2180 ( .A1(\RegFilePlugin_regFile[2][27] ), .A2(n1628), .B1(
        \RegFilePlugin_regFile[29][27] ), .B2(n1501), .ZN(n1404) );
  aoi22d1 U2181 ( .A1(\RegFilePlugin_regFile[16][27] ), .A2(n1975), .B1(
        \RegFilePlugin_regFile[17][27] ), .B2(n1953), .ZN(n1411) );
  aoi22d1 U2182 ( .A1(\RegFilePlugin_regFile[0][27] ), .A2(n2030), .B1(
        \RegFilePlugin_regFile[15][27] ), .B2(n2023), .ZN(n1410) );
  aoi22d1 U2183 ( .A1(\RegFilePlugin_regFile[26][27] ), .A2(n1649), .B1(
        \RegFilePlugin_regFile[8][27] ), .B2(n1902), .ZN(n1409) );
  aoi22d1 U2184 ( .A1(\RegFilePlugin_regFile[10][27] ), .A2(n1993), .B1(
        \RegFilePlugin_regFile[23][27] ), .B2(n2021), .ZN(n1408) );
  or04d0 U2185 ( .A1(n1415), .A2(n1414), .A3(n1413), .A4(n1412), .Z(N860) );
  aoi22d1 U2186 ( .A1(\RegFilePlugin_regFile[10][26] ), .A2(n1416), .B1(
        \RegFilePlugin_regFile[3][26] ), .B2(n1816), .ZN(n1421) );
  aoi22d1 U2187 ( .A1(\RegFilePlugin_regFile[29][26] ), .A2(n1974), .B1(
        \RegFilePlugin_regFile[16][26] ), .B2(n1671), .ZN(n1420) );
  aoi22d1 U2188 ( .A1(\RegFilePlugin_regFile[9][26] ), .A2(n1858), .B1(
        \RegFilePlugin_regFile[20][26] ), .B2(n2006), .ZN(n1419) );
  aoi22d1 U2189 ( .A1(\RegFilePlugin_regFile[31][26] ), .A2(n1417), .B1(
        \RegFilePlugin_regFile[21][26] ), .B2(n1931), .ZN(n1418) );
  aoi22d1 U2190 ( .A1(\RegFilePlugin_regFile[22][26] ), .A2(n1472), .B1(
        \RegFilePlugin_regFile[18][26] ), .B2(n1937), .ZN(n1425) );
  aoi22d1 U2191 ( .A1(\RegFilePlugin_regFile[8][26] ), .A2(n1670), .B1(
        \RegFilePlugin_regFile[27][26] ), .B2(n1718), .ZN(n1424) );
  aoi22d1 U2192 ( .A1(\RegFilePlugin_regFile[26][26] ), .A2(n2015), .B1(
        \RegFilePlugin_regFile[13][26] ), .B2(n2025), .ZN(n1423) );
  aoi22d1 U2193 ( .A1(\RegFilePlugin_regFile[6][26] ), .A2(n1522), .B1(
        \RegFilePlugin_regFile[7][26] ), .B2(n1925), .ZN(n1422) );
  aoi22d1 U2194 ( .A1(\RegFilePlugin_regFile[15][26] ), .A2(n1994), .B1(
        \RegFilePlugin_regFile[1][26] ), .B2(n2012), .ZN(n1429) );
  aoi22d1 U2195 ( .A1(\RegFilePlugin_regFile[25][26] ), .A2(n1926), .B1(
        \RegFilePlugin_regFile[11][26] ), .B2(n2013), .ZN(n1428) );
  aoi22d1 U2196 ( .A1(\RegFilePlugin_regFile[23][26] ), .A2(n1544), .B1(
        \RegFilePlugin_regFile[2][26] ), .B2(n1628), .ZN(n1427) );
  aoi22d1 U2197 ( .A1(\RegFilePlugin_regFile[5][26] ), .A2(n1606), .B1(
        \RegFilePlugin_regFile[28][26] ), .B2(n1892), .ZN(n1426) );
  aoi22d1 U2198 ( .A1(\RegFilePlugin_regFile[19][26] ), .A2(n2024), .B1(
        \RegFilePlugin_regFile[24][26] ), .B2(n2020), .ZN(n1433) );
  aoi22d1 U2199 ( .A1(\RegFilePlugin_regFile[17][26] ), .A2(n1953), .B1(
        \RegFilePlugin_regFile[4][26] ), .B2(n2004), .ZN(n1432) );
  aoi22d1 U2200 ( .A1(\RegFilePlugin_regFile[14][26] ), .A2(n1916), .B1(
        \RegFilePlugin_regFile[12][26] ), .B2(n2031), .ZN(n1431) );
  aoi22d1 U2201 ( .A1(\RegFilePlugin_regFile[30][26] ), .A2(n1987), .B1(
        \RegFilePlugin_regFile[0][26] ), .B2(n1585), .ZN(n1430) );
  or04d0 U2202 ( .A1(n1437), .A2(n1436), .A3(n1435), .A4(n1434), .Z(N861) );
  aoi22d1 U2203 ( .A1(\RegFilePlugin_regFile[14][29] ), .A2(n2003), .B1(
        \RegFilePlugin_regFile[20][29] ), .B2(n2006), .ZN(n1441) );
  aoi22d1 U2204 ( .A1(\RegFilePlugin_regFile[2][29] ), .A2(n2032), .B1(
        \RegFilePlugin_regFile[23][29] ), .B2(n1544), .ZN(n1440) );
  aoi22d1 U2205 ( .A1(\RegFilePlugin_regFile[13][29] ), .A2(n1932), .B1(
        \RegFilePlugin_regFile[3][29] ), .B2(n2022), .ZN(n1439) );
  aoi22d1 U2206 ( .A1(\RegFilePlugin_regFile[5][29] ), .A2(n1606), .B1(
        \RegFilePlugin_regFile[10][29] ), .B2(n1993), .ZN(n1438) );
  aoi22d1 U2207 ( .A1(\RegFilePlugin_regFile[9][29] ), .A2(n2011), .B1(
        \RegFilePlugin_regFile[8][29] ), .B2(n1670), .ZN(n1445) );
  aoi22d1 U2208 ( .A1(\RegFilePlugin_regFile[21][29] ), .A2(n1931), .B1(
        \RegFilePlugin_regFile[30][29] ), .B2(n1987), .ZN(n1444) );
  aoi22d1 U2209 ( .A1(\RegFilePlugin_regFile[27][29] ), .A2(n2033), .B1(
        \RegFilePlugin_regFile[17][29] ), .B2(n1953), .ZN(n1443) );
  aoi22d1 U2210 ( .A1(\RegFilePlugin_regFile[18][29] ), .A2(n1937), .B1(
        \RegFilePlugin_regFile[26][29] ), .B2(n1649), .ZN(n1442) );
  aoi22d1 U2211 ( .A1(\RegFilePlugin_regFile[31][29] ), .A2(n1942), .B1(
        \RegFilePlugin_regFile[29][29] ), .B2(n1501), .ZN(n1449) );
  aoi22d1 U2212 ( .A1(\RegFilePlugin_regFile[15][29] ), .A2(n2023), .B1(
        \RegFilePlugin_regFile[12][29] ), .B2(n2031), .ZN(n1448) );
  aoi22d1 U2213 ( .A1(\RegFilePlugin_regFile[1][29] ), .A2(n1692), .B1(
        \RegFilePlugin_regFile[6][29] ), .B2(n1943), .ZN(n1447) );
  aoi22d1 U2214 ( .A1(\RegFilePlugin_regFile[16][29] ), .A2(n1975), .B1(
        \RegFilePlugin_regFile[7][29] ), .B2(n1925), .ZN(n1446) );
  aoi22d1 U2215 ( .A1(\RegFilePlugin_regFile[0][29] ), .A2(n2030), .B1(
        \RegFilePlugin_regFile[11][29] ), .B2(n2013), .ZN(n1453) );
  aoi22d1 U2216 ( .A1(\RegFilePlugin_regFile[24][29] ), .A2(n2020), .B1(
        \RegFilePlugin_regFile[4][29] ), .B2(n2004), .ZN(n1452) );
  aoi22d1 U2217 ( .A1(\RegFilePlugin_regFile[22][29] ), .A2(n2014), .B1(
        \RegFilePlugin_regFile[19][29] ), .B2(n2024), .ZN(n1451) );
  aoi22d1 U2218 ( .A1(\RegFilePlugin_regFile[25][29] ), .A2(n1926), .B1(
        \RegFilePlugin_regFile[28][29] ), .B2(n1892), .ZN(n1450) );
  or04d0 U2219 ( .A1(n1457), .A2(n1456), .A3(n1455), .A4(n1454), .Z(N858) );
  aoi22d1 U2220 ( .A1(\RegFilePlugin_regFile[2][19] ), .A2(n2032), .B1(
        \RegFilePlugin_regFile[21][19] ), .B2(n1377), .ZN(n1462) );
  aoi22d1 U2221 ( .A1(\RegFilePlugin_regFile[31][19] ), .A2(n1942), .B1(
        \RegFilePlugin_regFile[14][19] ), .B2(n1916), .ZN(n1461) );
  aoi22d1 U2222 ( .A1(\RegFilePlugin_regFile[1][19] ), .A2(n2012), .B1(
        \RegFilePlugin_regFile[27][19] ), .B2(n1718), .ZN(n1460) );
  aoi22d1 U2223 ( .A1(\RegFilePlugin_regFile[7][19] ), .A2(n1925), .B1(
        \RegFilePlugin_regFile[19][19] ), .B2(n1458), .ZN(n1459) );
  aoi22d1 U2224 ( .A1(\RegFilePlugin_regFile[25][19] ), .A2(n1926), .B1(
        \RegFilePlugin_regFile[28][19] ), .B2(n1903), .ZN(n1467) );
  aoi22d1 U2225 ( .A1(\RegFilePlugin_regFile[9][19] ), .A2(n1858), .B1(
        \RegFilePlugin_regFile[6][19] ), .B2(n1943), .ZN(n1466) );
  buffd1 U2226 ( .I(n1463), .Z(n1981) );
  aoi22d1 U2227 ( .A1(\RegFilePlugin_regFile[12][19] ), .A2(n1981), .B1(
        \RegFilePlugin_regFile[10][19] ), .B2(n1416), .ZN(n1465) );
  aoi22d1 U2228 ( .A1(\RegFilePlugin_regFile[0][19] ), .A2(n2030), .B1(
        \RegFilePlugin_regFile[3][19] ), .B2(n1816), .ZN(n1464) );
  aoi22d1 U2229 ( .A1(\RegFilePlugin_regFile[30][19] ), .A2(n1987), .B1(
        \RegFilePlugin_regFile[17][19] ), .B2(n1953), .ZN(n1471) );
  aoi22d1 U2230 ( .A1(\RegFilePlugin_regFile[23][19] ), .A2(n2021), .B1(
        \RegFilePlugin_regFile[29][19] ), .B2(n1974), .ZN(n1470) );
  aoi22d1 U2231 ( .A1(\RegFilePlugin_regFile[11][19] ), .A2(n2013), .B1(
        \RegFilePlugin_regFile[16][19] ), .B2(n1671), .ZN(n1469) );
  aoi22d1 U2232 ( .A1(\RegFilePlugin_regFile[18][19] ), .A2(n1937), .B1(
        \RegFilePlugin_regFile[24][19] ), .B2(n2020), .ZN(n1468) );
  aoi22d1 U2233 ( .A1(\RegFilePlugin_regFile[5][19] ), .A2(n1982), .B1(
        \RegFilePlugin_regFile[4][19] ), .B2(n1879), .ZN(n1476) );
  aoi22d1 U2234 ( .A1(\RegFilePlugin_regFile[15][19] ), .A2(n2023), .B1(
        \RegFilePlugin_regFile[26][19] ), .B2(n1649), .ZN(n1475) );
  aoi22d1 U2235 ( .A1(\RegFilePlugin_regFile[20][19] ), .A2(n2006), .B1(
        \RegFilePlugin_regFile[8][19] ), .B2(n1670), .ZN(n1474) );
  buffd1 U2236 ( .I(n1472), .Z(n1988) );
  aoi22d1 U2237 ( .A1(\RegFilePlugin_regFile[13][19] ), .A2(n2025), .B1(
        \RegFilePlugin_regFile[22][19] ), .B2(n1988), .ZN(n1473) );
  or04d0 U2238 ( .A1(n1480), .A2(n1479), .A3(n1478), .A4(n1477), .Z(N868) );
  aoi22d1 U2239 ( .A1(\RegFilePlugin_regFile[20][23] ), .A2(n1387), .B1(
        \RegFilePlugin_regFile[18][23] ), .B2(n1937), .ZN(n1484) );
  aoi22d1 U2240 ( .A1(\RegFilePlugin_regFile[22][23] ), .A2(n1988), .B1(
        \RegFilePlugin_regFile[24][23] ), .B2(n2020), .ZN(n1483) );
  aoi22d1 U2241 ( .A1(\RegFilePlugin_regFile[10][23] ), .A2(n1416), .B1(
        \RegFilePlugin_regFile[21][23] ), .B2(n1931), .ZN(n1482) );
  aoi22d1 U2242 ( .A1(\RegFilePlugin_regFile[23][23] ), .A2(n1544), .B1(
        \RegFilePlugin_regFile[31][23] ), .B2(n1942), .ZN(n1481) );
  aoi22d1 U2243 ( .A1(\RegFilePlugin_regFile[26][23] ), .A2(n2015), .B1(
        \RegFilePlugin_regFile[13][23] ), .B2(n1932), .ZN(n1488) );
  aoi22d1 U2244 ( .A1(\RegFilePlugin_regFile[4][23] ), .A2(n2004), .B1(
        \RegFilePlugin_regFile[30][23] ), .B2(n1837), .ZN(n1487) );
  aoi22d1 U2245 ( .A1(\RegFilePlugin_regFile[16][23] ), .A2(n1975), .B1(
        \RegFilePlugin_regFile[9][23] ), .B2(n2011), .ZN(n1486) );
  aoi22d1 U2246 ( .A1(\RegFilePlugin_regFile[2][23] ), .A2(n2032), .B1(
        \RegFilePlugin_regFile[6][23] ), .B2(n1943), .ZN(n1485) );
  aoi22d1 U2247 ( .A1(\RegFilePlugin_regFile[7][23] ), .A2(n1543), .B1(
        \RegFilePlugin_regFile[11][23] ), .B2(n2013), .ZN(n1492) );
  aoi22d1 U2248 ( .A1(\RegFilePlugin_regFile[27][23] ), .A2(n1718), .B1(
        \RegFilePlugin_regFile[8][23] ), .B2(n1902), .ZN(n1491) );
  aoi22d1 U2249 ( .A1(\RegFilePlugin_regFile[0][23] ), .A2(n2030), .B1(
        \RegFilePlugin_regFile[17][23] ), .B2(n1953), .ZN(n1490) );
  aoi22d1 U2250 ( .A1(\RegFilePlugin_regFile[19][23] ), .A2(n2024), .B1(
        \RegFilePlugin_regFile[28][23] ), .B2(n1892), .ZN(n1489) );
  aoi22d1 U2251 ( .A1(\RegFilePlugin_regFile[25][23] ), .A2(n1607), .B1(
        \RegFilePlugin_regFile[12][23] ), .B2(n1981), .ZN(n1496) );
  aoi22d1 U2252 ( .A1(\RegFilePlugin_regFile[3][23] ), .A2(n1816), .B1(
        \RegFilePlugin_regFile[29][23] ), .B2(n1501), .ZN(n1495) );
  aoi22d1 U2253 ( .A1(\RegFilePlugin_regFile[14][23] ), .A2(n1916), .B1(
        \RegFilePlugin_regFile[1][23] ), .B2(n2012), .ZN(n1494) );
  aoi22d1 U2254 ( .A1(\RegFilePlugin_regFile[15][23] ), .A2(n2023), .B1(
        \RegFilePlugin_regFile[5][23] ), .B2(n1982), .ZN(n1493) );
  or04d0 U2255 ( .A1(n1500), .A2(n1499), .A3(n1498), .A4(n1497), .Z(N864) );
  aoi22d1 U2256 ( .A1(\RegFilePlugin_regFile[29][6] ), .A2(n1501), .B1(
        \RegFilePlugin_regFile[16][6] ), .B2(n1975), .ZN(n1505) );
  aoi22d1 U2257 ( .A1(\RegFilePlugin_regFile[30][6] ), .A2(n1837), .B1(
        \RegFilePlugin_regFile[18][6] ), .B2(n1952), .ZN(n1504) );
  aoi22d1 U2258 ( .A1(\RegFilePlugin_regFile[26][6] ), .A2(n2015), .B1(
        \RegFilePlugin_regFile[4][6] ), .B2(n2004), .ZN(n1503) );
  aoi22d1 U2259 ( .A1(\RegFilePlugin_regFile[9][6] ), .A2(n1858), .B1(
        \RegFilePlugin_regFile[31][6] ), .B2(n1942), .ZN(n1502) );
  aoi22d1 U2260 ( .A1(\RegFilePlugin_regFile[12][6] ), .A2(n2031), .B1(
        \RegFilePlugin_regFile[6][6] ), .B2(n1943), .ZN(n1509) );
  aoi22d1 U2261 ( .A1(\RegFilePlugin_regFile[23][6] ), .A2(n2021), .B1(
        \RegFilePlugin_regFile[20][6] ), .B2(n2006), .ZN(n1508) );
  aoi22d1 U2262 ( .A1(\RegFilePlugin_regFile[25][6] ), .A2(n1926), .B1(
        \RegFilePlugin_regFile[7][6] ), .B2(n1925), .ZN(n1507) );
  aoi22d1 U2263 ( .A1(\RegFilePlugin_regFile[28][6] ), .A2(n1903), .B1(
        \RegFilePlugin_regFile[22][6] ), .B2(n1988), .ZN(n1506) );
  aoi22d1 U2264 ( .A1(\RegFilePlugin_regFile[1][6] ), .A2(n2012), .B1(
        \RegFilePlugin_regFile[3][6] ), .B2(n2022), .ZN(n1513) );
  aoi22d1 U2265 ( .A1(\RegFilePlugin_regFile[14][6] ), .A2(n2003), .B1(
        \RegFilePlugin_regFile[13][6] ), .B2(n2025), .ZN(n1512) );
  aoi22d1 U2266 ( .A1(\RegFilePlugin_regFile[17][6] ), .A2(n1953), .B1(
        \RegFilePlugin_regFile[8][6] ), .B2(n1670), .ZN(n1511) );
  aoi22d1 U2267 ( .A1(\RegFilePlugin_regFile[2][6] ), .A2(n2032), .B1(
        \RegFilePlugin_regFile[5][6] ), .B2(n1982), .ZN(n1510) );
  aoi22d1 U2268 ( .A1(\RegFilePlugin_regFile[15][6] ), .A2(n1994), .B1(
        \RegFilePlugin_regFile[10][6] ), .B2(n1993), .ZN(n1517) );
  aoi22d1 U2269 ( .A1(\RegFilePlugin_regFile[11][6] ), .A2(n2013), .B1(
        \RegFilePlugin_regFile[24][6] ), .B2(n1735), .ZN(n1516) );
  aoi22d1 U2270 ( .A1(\RegFilePlugin_regFile[19][6] ), .A2(n2024), .B1(
        \RegFilePlugin_regFile[27][6] ), .B2(n2033), .ZN(n1515) );
  aoi22d1 U2271 ( .A1(\RegFilePlugin_regFile[0][6] ), .A2(n2030), .B1(
        \RegFilePlugin_regFile[21][6] ), .B2(n1931), .ZN(n1514) );
  or04d0 U2272 ( .A1(n1521), .A2(n1520), .A3(n1519), .A4(n1518), .Z(N881) );
  aoi22d1 U2273 ( .A1(\RegFilePlugin_regFile[26][21] ), .A2(n1649), .B1(
        \RegFilePlugin_regFile[29][21] ), .B2(n1974), .ZN(n1526) );
  aoi22d1 U2274 ( .A1(\RegFilePlugin_regFile[17][21] ), .A2(n1976), .B1(
        \RegFilePlugin_regFile[6][21] ), .B2(n1522), .ZN(n1525) );
  aoi22d1 U2275 ( .A1(\RegFilePlugin_regFile[0][21] ), .A2(n2030), .B1(
        \RegFilePlugin_regFile[25][21] ), .B2(n1607), .ZN(n1524) );
  aoi22d1 U2276 ( .A1(\RegFilePlugin_regFile[12][21] ), .A2(n1981), .B1(
        \RegFilePlugin_regFile[16][21] ), .B2(n1671), .ZN(n1523) );
  aoi22d1 U2277 ( .A1(\RegFilePlugin_regFile[24][21] ), .A2(n1735), .B1(
        \RegFilePlugin_regFile[7][21] ), .B2(n1925), .ZN(n1530) );
  aoi22d1 U2278 ( .A1(\RegFilePlugin_regFile[3][21] ), .A2(n1816), .B1(
        \RegFilePlugin_regFile[4][21] ), .B2(n1879), .ZN(n1529) );
  aoi22d1 U2279 ( .A1(\RegFilePlugin_regFile[23][21] ), .A2(n2021), .B1(
        \RegFilePlugin_regFile[9][21] ), .B2(n1858), .ZN(n1528) );
  aoi22d1 U2280 ( .A1(\RegFilePlugin_regFile[15][21] ), .A2(n2023), .B1(
        \RegFilePlugin_regFile[28][21] ), .B2(n1892), .ZN(n1527) );
  aoi22d1 U2281 ( .A1(\RegFilePlugin_regFile[20][21] ), .A2(n1387), .B1(
        \RegFilePlugin_regFile[11][21] ), .B2(n2013), .ZN(n1534) );
  aoi22d1 U2282 ( .A1(\RegFilePlugin_regFile[2][21] ), .A2(n2032), .B1(
        \RegFilePlugin_regFile[5][21] ), .B2(n1982), .ZN(n1533) );
  aoi22d1 U2283 ( .A1(\RegFilePlugin_regFile[31][21] ), .A2(n1942), .B1(
        \RegFilePlugin_regFile[30][21] ), .B2(n1837), .ZN(n1532) );
  aoi22d1 U2284 ( .A1(\RegFilePlugin_regFile[27][21] ), .A2(n2033), .B1(
        \RegFilePlugin_regFile[18][21] ), .B2(n1937), .ZN(n1531) );
  aoi22d1 U2285 ( .A1(\RegFilePlugin_regFile[13][21] ), .A2(n1932), .B1(
        \RegFilePlugin_regFile[21][21] ), .B2(n1377), .ZN(n1538) );
  aoi22d1 U2286 ( .A1(\RegFilePlugin_regFile[8][21] ), .A2(n1902), .B1(
        \RegFilePlugin_regFile[22][21] ), .B2(n1988), .ZN(n1537) );
  aoi22d1 U2287 ( .A1(\RegFilePlugin_regFile[10][21] ), .A2(n1993), .B1(
        \RegFilePlugin_regFile[19][21] ), .B2(n1458), .ZN(n1536) );
  aoi22d1 U2288 ( .A1(\RegFilePlugin_regFile[14][21] ), .A2(n1916), .B1(
        \RegFilePlugin_regFile[1][21] ), .B2(n1692), .ZN(n1535) );
  or04d0 U2289 ( .A1(n1542), .A2(n1541), .A3(n1540), .A4(n1539), .Z(N866) );
  aoi22d1 U2290 ( .A1(\RegFilePlugin_regFile[12][15] ), .A2(n1981), .B1(
        \RegFilePlugin_regFile[30][15] ), .B2(n1837), .ZN(n1548) );
  aoi22d1 U2291 ( .A1(\RegFilePlugin_regFile[8][15] ), .A2(n1670), .B1(
        \RegFilePlugin_regFile[7][15] ), .B2(n1543), .ZN(n1547) );
  aoi22d1 U2292 ( .A1(\RegFilePlugin_regFile[23][15] ), .A2(n1544), .B1(
        \RegFilePlugin_regFile[4][15] ), .B2(n2004), .ZN(n1546) );
  aoi22d1 U2293 ( .A1(\RegFilePlugin_regFile[27][15] ), .A2(n2033), .B1(
        \RegFilePlugin_regFile[25][15] ), .B2(n1607), .ZN(n1545) );
  aoi22d1 U2294 ( .A1(\RegFilePlugin_regFile[16][15] ), .A2(n1671), .B1(
        \RegFilePlugin_regFile[18][15] ), .B2(n1937), .ZN(n1552) );
  aoi22d1 U2295 ( .A1(\RegFilePlugin_regFile[24][15] ), .A2(n1735), .B1(
        \RegFilePlugin_regFile[10][15] ), .B2(n1416), .ZN(n1551) );
  aoi22d1 U2296 ( .A1(\RegFilePlugin_regFile[2][15] ), .A2(n2032), .B1(
        \RegFilePlugin_regFile[5][15] ), .B2(n1606), .ZN(n1550) );
  aoi22d1 U2297 ( .A1(\RegFilePlugin_regFile[11][15] ), .A2(n1901), .B1(
        \RegFilePlugin_regFile[9][15] ), .B2(n1858), .ZN(n1549) );
  aoi22d1 U2298 ( .A1(\RegFilePlugin_regFile[26][15] ), .A2(n2015), .B1(
        \RegFilePlugin_regFile[22][15] ), .B2(n1988), .ZN(n1556) );
  aoi22d1 U2299 ( .A1(\RegFilePlugin_regFile[3][15] ), .A2(n1816), .B1(
        \RegFilePlugin_regFile[1][15] ), .B2(n1692), .ZN(n1555) );
  aoi22d1 U2300 ( .A1(\RegFilePlugin_regFile[29][15] ), .A2(n1501), .B1(
        \RegFilePlugin_regFile[14][15] ), .B2(n1916), .ZN(n1554) );
  aoi22d1 U2301 ( .A1(\RegFilePlugin_regFile[31][15] ), .A2(n1417), .B1(
        \RegFilePlugin_regFile[17][15] ), .B2(n1953), .ZN(n1553) );
  aoi22d1 U2302 ( .A1(\RegFilePlugin_regFile[19][15] ), .A2(n2024), .B1(
        \RegFilePlugin_regFile[21][15] ), .B2(n1377), .ZN(n1560) );
  aoi22d1 U2303 ( .A1(\RegFilePlugin_regFile[15][15] ), .A2(n2023), .B1(
        \RegFilePlugin_regFile[28][15] ), .B2(n1892), .ZN(n1559) );
  aoi22d1 U2304 ( .A1(\RegFilePlugin_regFile[13][15] ), .A2(n2025), .B1(
        \RegFilePlugin_regFile[0][15] ), .B2(n1585), .ZN(n1558) );
  aoi22d1 U2305 ( .A1(\RegFilePlugin_regFile[6][15] ), .A2(n1522), .B1(
        \RegFilePlugin_regFile[20][15] ), .B2(n2006), .ZN(n1557) );
  or04d0 U2306 ( .A1(n1564), .A2(n1563), .A3(n1562), .A4(n1561), .Z(N872) );
  aoi22d1 U2307 ( .A1(\RegFilePlugin_regFile[1][30] ), .A2(n2012), .B1(
        \RegFilePlugin_regFile[12][30] ), .B2(n2031), .ZN(n1568) );
  aoi22d1 U2308 ( .A1(\RegFilePlugin_regFile[21][30] ), .A2(n1931), .B1(
        \RegFilePlugin_regFile[20][30] ), .B2(n1387), .ZN(n1567) );
  aoi22d1 U2309 ( .A1(\RegFilePlugin_regFile[13][30] ), .A2(n2025), .B1(
        \RegFilePlugin_regFile[19][30] ), .B2(n2024), .ZN(n1566) );
  aoi22d1 U2310 ( .A1(\RegFilePlugin_regFile[16][30] ), .A2(n1671), .B1(
        \RegFilePlugin_regFile[4][30] ), .B2(n1879), .ZN(n1565) );
  aoi22d1 U2311 ( .A1(\RegFilePlugin_regFile[27][30] ), .A2(n2033), .B1(
        \RegFilePlugin_regFile[7][30] ), .B2(n1543), .ZN(n1572) );
  aoi22d1 U2312 ( .A1(\RegFilePlugin_regFile[8][30] ), .A2(n1902), .B1(
        \RegFilePlugin_regFile[17][30] ), .B2(n1976), .ZN(n1571) );
  aoi22d1 U2313 ( .A1(\RegFilePlugin_regFile[5][30] ), .A2(n1982), .B1(
        \RegFilePlugin_regFile[2][30] ), .B2(n1628), .ZN(n1570) );
  aoi22d1 U2314 ( .A1(\RegFilePlugin_regFile[30][30] ), .A2(n1837), .B1(
        \RegFilePlugin_regFile[15][30] ), .B2(n2023), .ZN(n1569) );
  aoi22d1 U2315 ( .A1(\RegFilePlugin_regFile[25][30] ), .A2(n1926), .B1(
        \RegFilePlugin_regFile[0][30] ), .B2(n1585), .ZN(n1576) );
  aoi22d1 U2316 ( .A1(\RegFilePlugin_regFile[10][30] ), .A2(n1993), .B1(
        \RegFilePlugin_regFile[11][30] ), .B2(n2013), .ZN(n1575) );
  aoi22d1 U2317 ( .A1(\RegFilePlugin_regFile[3][30] ), .A2(n1816), .B1(
        \RegFilePlugin_regFile[29][30] ), .B2(n1501), .ZN(n1574) );
  aoi22d1 U2318 ( .A1(\RegFilePlugin_regFile[14][30] ), .A2(n1916), .B1(
        \RegFilePlugin_regFile[31][30] ), .B2(n1942), .ZN(n1573) );
  aoi22d1 U2319 ( .A1(\RegFilePlugin_regFile[6][30] ), .A2(n1522), .B1(
        \RegFilePlugin_regFile[26][30] ), .B2(n2015), .ZN(n1580) );
  aoi22d1 U2320 ( .A1(\RegFilePlugin_regFile[23][30] ), .A2(n2021), .B1(
        \RegFilePlugin_regFile[22][30] ), .B2(n2014), .ZN(n1579) );
  aoi22d1 U2321 ( .A1(\RegFilePlugin_regFile[24][30] ), .A2(n2020), .B1(
        \RegFilePlugin_regFile[9][30] ), .B2(n2011), .ZN(n1578) );
  aoi22d1 U2322 ( .A1(\RegFilePlugin_regFile[18][30] ), .A2(n1937), .B1(
        \RegFilePlugin_regFile[28][30] ), .B2(n1903), .ZN(n1577) );
  or04d0 U2323 ( .A1(n1584), .A2(n1583), .A3(n1582), .A4(n1581), .Z(N857) );
  aoi22d1 U2324 ( .A1(\RegFilePlugin_regFile[7][20] ), .A2(n1925), .B1(
        \RegFilePlugin_regFile[4][20] ), .B2(n1879), .ZN(n1589) );
  aoi22d1 U2325 ( .A1(\RegFilePlugin_regFile[23][20] ), .A2(n2021), .B1(
        \RegFilePlugin_regFile[0][20] ), .B2(n1585), .ZN(n1588) );
  aoi22d1 U2326 ( .A1(\RegFilePlugin_regFile[3][20] ), .A2(n2022), .B1(
        \RegFilePlugin_regFile[10][20] ), .B2(n1416), .ZN(n1587) );
  aoi22d1 U2327 ( .A1(\RegFilePlugin_regFile[19][20] ), .A2(n2024), .B1(
        \RegFilePlugin_regFile[5][20] ), .B2(n1982), .ZN(n1586) );
  aoi22d1 U2328 ( .A1(\RegFilePlugin_regFile[20][20] ), .A2(n1387), .B1(
        \RegFilePlugin_regFile[22][20] ), .B2(n1988), .ZN(n1593) );
  aoi22d1 U2329 ( .A1(\RegFilePlugin_regFile[13][20] ), .A2(n2025), .B1(
        \RegFilePlugin_regFile[29][20] ), .B2(n1974), .ZN(n1592) );
  aoi22d1 U2330 ( .A1(\RegFilePlugin_regFile[24][20] ), .A2(n1735), .B1(
        \RegFilePlugin_regFile[27][20] ), .B2(n1718), .ZN(n1591) );
  aoi22d1 U2331 ( .A1(\RegFilePlugin_regFile[9][20] ), .A2(n2011), .B1(
        \RegFilePlugin_regFile[18][20] ), .B2(n1952), .ZN(n1590) );
  aoi22d1 U2332 ( .A1(\RegFilePlugin_regFile[30][20] ), .A2(n1987), .B1(
        \RegFilePlugin_regFile[17][20] ), .B2(n1953), .ZN(n1597) );
  aoi22d1 U2333 ( .A1(\RegFilePlugin_regFile[2][20] ), .A2(n2032), .B1(
        \RegFilePlugin_regFile[21][20] ), .B2(n1931), .ZN(n1596) );
  aoi22d1 U2334 ( .A1(\RegFilePlugin_regFile[28][20] ), .A2(n1892), .B1(
        \RegFilePlugin_regFile[6][20] ), .B2(n1943), .ZN(n1595) );
  aoi22d1 U2335 ( .A1(\RegFilePlugin_regFile[31][20] ), .A2(n1942), .B1(
        \RegFilePlugin_regFile[11][20] ), .B2(n2013), .ZN(n1594) );
  aoi22d1 U2336 ( .A1(\RegFilePlugin_regFile[14][20] ), .A2(n2003), .B1(
        \RegFilePlugin_regFile[12][20] ), .B2(n1981), .ZN(n1601) );
  aoi22d1 U2337 ( .A1(\RegFilePlugin_regFile[25][20] ), .A2(n1926), .B1(
        \RegFilePlugin_regFile[8][20] ), .B2(n1902), .ZN(n1600) );
  aoi22d1 U2338 ( .A1(\RegFilePlugin_regFile[26][20] ), .A2(n1649), .B1(
        \RegFilePlugin_regFile[15][20] ), .B2(n1994), .ZN(n1599) );
  aoi22d1 U2339 ( .A1(\RegFilePlugin_regFile[1][20] ), .A2(n2012), .B1(
        \RegFilePlugin_regFile[16][20] ), .B2(n1671), .ZN(n1598) );
  or04d0 U2340 ( .A1(n1605), .A2(n1604), .A3(n1603), .A4(n1602), .Z(N867) );
  aoi22d1 U2341 ( .A1(\RegFilePlugin_regFile[4][25] ), .A2(n2004), .B1(
        \RegFilePlugin_regFile[9][25] ), .B2(n2011), .ZN(n1611) );
  aoi22d1 U2342 ( .A1(\RegFilePlugin_regFile[16][25] ), .A2(n1671), .B1(
        \RegFilePlugin_regFile[5][25] ), .B2(n1606), .ZN(n1610) );
  aoi22d1 U2343 ( .A1(\RegFilePlugin_regFile[23][25] ), .A2(n1544), .B1(
        \RegFilePlugin_regFile[6][25] ), .B2(n1522), .ZN(n1609) );
  aoi22d1 U2344 ( .A1(\RegFilePlugin_regFile[25][25] ), .A2(n1607), .B1(
        \RegFilePlugin_regFile[8][25] ), .B2(n1902), .ZN(n1608) );
  aoi22d1 U2345 ( .A1(\RegFilePlugin_regFile[0][25] ), .A2(n2030), .B1(
        \RegFilePlugin_regFile[2][25] ), .B2(n1628), .ZN(n1615) );
  aoi22d1 U2346 ( .A1(\RegFilePlugin_regFile[31][25] ), .A2(n1417), .B1(
        \RegFilePlugin_regFile[10][25] ), .B2(n1416), .ZN(n1614) );
  aoi22d1 U2347 ( .A1(\RegFilePlugin_regFile[28][25] ), .A2(n1892), .B1(
        \RegFilePlugin_regFile[27][25] ), .B2(n1718), .ZN(n1613) );
  aoi22d1 U2348 ( .A1(\RegFilePlugin_regFile[30][25] ), .A2(n1987), .B1(
        \RegFilePlugin_regFile[18][25] ), .B2(n1937), .ZN(n1612) );
  aoi22d1 U2349 ( .A1(\RegFilePlugin_regFile[3][25] ), .A2(n1816), .B1(
        \RegFilePlugin_regFile[12][25] ), .B2(n2031), .ZN(n1619) );
  aoi22d1 U2350 ( .A1(\RegFilePlugin_regFile[7][25] ), .A2(n1543), .B1(
        \RegFilePlugin_regFile[19][25] ), .B2(n1458), .ZN(n1618) );
  aoi22d1 U2351 ( .A1(\RegFilePlugin_regFile[17][25] ), .A2(n1976), .B1(
        \RegFilePlugin_regFile[13][25] ), .B2(n1932), .ZN(n1617) );
  aoi22d1 U2352 ( .A1(\RegFilePlugin_regFile[29][25] ), .A2(n1974), .B1(
        \RegFilePlugin_regFile[15][25] ), .B2(n2023), .ZN(n1616) );
  aoi22d1 U2353 ( .A1(\RegFilePlugin_regFile[20][25] ), .A2(n1387), .B1(
        \RegFilePlugin_regFile[11][25] ), .B2(n2013), .ZN(n1623) );
  aoi22d1 U2354 ( .A1(\RegFilePlugin_regFile[21][25] ), .A2(n1377), .B1(
        \RegFilePlugin_regFile[1][25] ), .B2(n1692), .ZN(n1622) );
  aoi22d1 U2355 ( .A1(\RegFilePlugin_regFile[14][25] ), .A2(n2003), .B1(
        \RegFilePlugin_regFile[22][25] ), .B2(n2014), .ZN(n1621) );
  aoi22d1 U2356 ( .A1(\RegFilePlugin_regFile[26][25] ), .A2(n1649), .B1(
        \RegFilePlugin_regFile[24][25] ), .B2(n2020), .ZN(n1620) );
  or04d0 U2357 ( .A1(n1627), .A2(n1626), .A3(n1625), .A4(n1624), .Z(N862) );
  aoi22d1 U2358 ( .A1(\RegFilePlugin_regFile[14][5] ), .A2(n2003), .B1(
        \RegFilePlugin_regFile[2][5] ), .B2(n1628), .ZN(n1632) );
  aoi22d1 U2359 ( .A1(\RegFilePlugin_regFile[15][5] ), .A2(n1994), .B1(
        \RegFilePlugin_regFile[17][5] ), .B2(n1976), .ZN(n1631) );
  aoi22d1 U2360 ( .A1(\RegFilePlugin_regFile[8][5] ), .A2(n1902), .B1(
        \RegFilePlugin_regFile[26][5] ), .B2(n1649), .ZN(n1630) );
  aoi22d1 U2361 ( .A1(\RegFilePlugin_regFile[0][5] ), .A2(n2030), .B1(
        \RegFilePlugin_regFile[28][5] ), .B2(n1903), .ZN(n1629) );
  aoi22d1 U2362 ( .A1(\RegFilePlugin_regFile[22][5] ), .A2(n1988), .B1(
        \RegFilePlugin_regFile[19][5] ), .B2(n2024), .ZN(n1636) );
  aoi22d1 U2363 ( .A1(\RegFilePlugin_regFile[23][5] ), .A2(n1544), .B1(
        \RegFilePlugin_regFile[30][5] ), .B2(n1837), .ZN(n1635) );
  aoi22d1 U2364 ( .A1(\RegFilePlugin_regFile[16][5] ), .A2(n1671), .B1(
        \RegFilePlugin_regFile[31][5] ), .B2(n1417), .ZN(n1634) );
  aoi22d1 U2365 ( .A1(\RegFilePlugin_regFile[1][5] ), .A2(n1692), .B1(
        \RegFilePlugin_regFile[3][5] ), .B2(n2022), .ZN(n1633) );
  aoi22d1 U2366 ( .A1(\RegFilePlugin_regFile[11][5] ), .A2(n1901), .B1(
        \RegFilePlugin_regFile[18][5] ), .B2(n1952), .ZN(n1640) );
  aoi22d1 U2367 ( .A1(\RegFilePlugin_regFile[4][5] ), .A2(n2004), .B1(
        \RegFilePlugin_regFile[5][5] ), .B2(n1606), .ZN(n1639) );
  aoi22d1 U2368 ( .A1(\RegFilePlugin_regFile[12][5] ), .A2(n1981), .B1(
        \RegFilePlugin_regFile[7][5] ), .B2(n1925), .ZN(n1638) );
  aoi22d1 U2369 ( .A1(\RegFilePlugin_regFile[24][5] ), .A2(n2020), .B1(
        \RegFilePlugin_regFile[13][5] ), .B2(n2025), .ZN(n1637) );
  aoi22d1 U2370 ( .A1(\RegFilePlugin_regFile[6][5] ), .A2(n1522), .B1(
        \RegFilePlugin_regFile[10][5] ), .B2(n1993), .ZN(n1644) );
  aoi22d1 U2371 ( .A1(\RegFilePlugin_regFile[29][5] ), .A2(n1501), .B1(
        \RegFilePlugin_regFile[27][5] ), .B2(n2033), .ZN(n1643) );
  aoi22d1 U2372 ( .A1(\RegFilePlugin_regFile[9][5] ), .A2(n2011), .B1(
        \RegFilePlugin_regFile[25][5] ), .B2(n1607), .ZN(n1642) );
  aoi22d1 U2373 ( .A1(\RegFilePlugin_regFile[20][5] ), .A2(n1387), .B1(
        \RegFilePlugin_regFile[21][5] ), .B2(n1931), .ZN(n1641) );
  or04d0 U2374 ( .A1(n1648), .A2(n1647), .A3(n1646), .A4(n1645), .Z(N882) );
  aoi22d1 U2375 ( .A1(\RegFilePlugin_regFile[26][18] ), .A2(n1649), .B1(
        \RegFilePlugin_regFile[23][18] ), .B2(n2021), .ZN(n1653) );
  aoi22d1 U2376 ( .A1(\RegFilePlugin_regFile[4][18] ), .A2(n2004), .B1(
        \RegFilePlugin_regFile[6][18] ), .B2(n1943), .ZN(n1652) );
  aoi22d1 U2377 ( .A1(\RegFilePlugin_regFile[24][18] ), .A2(n1735), .B1(
        \RegFilePlugin_regFile[3][18] ), .B2(n2022), .ZN(n1651) );
  aoi22d1 U2378 ( .A1(\RegFilePlugin_regFile[22][18] ), .A2(n2014), .B1(
        \RegFilePlugin_regFile[18][18] ), .B2(n1952), .ZN(n1650) );
  aoi22d1 U2379 ( .A1(\RegFilePlugin_regFile[8][18] ), .A2(n1902), .B1(
        \RegFilePlugin_regFile[17][18] ), .B2(n1976), .ZN(n1657) );
  aoi22d1 U2380 ( .A1(\RegFilePlugin_regFile[11][18] ), .A2(n1901), .B1(
        \RegFilePlugin_regFile[31][18] ), .B2(n1942), .ZN(n1656) );
  aoi22d1 U2381 ( .A1(\RegFilePlugin_regFile[21][18] ), .A2(n1377), .B1(
        \RegFilePlugin_regFile[12][18] ), .B2(n1981), .ZN(n1655) );
  aoi22d1 U2382 ( .A1(\RegFilePlugin_regFile[16][18] ), .A2(n1975), .B1(
        \RegFilePlugin_regFile[14][18] ), .B2(n2003), .ZN(n1654) );
  aoi22d1 U2383 ( .A1(\RegFilePlugin_regFile[29][18] ), .A2(n1501), .B1(
        \RegFilePlugin_regFile[7][18] ), .B2(n1543), .ZN(n1661) );
  aoi22d1 U2384 ( .A1(\RegFilePlugin_regFile[1][18] ), .A2(n1692), .B1(
        \RegFilePlugin_regFile[28][18] ), .B2(n1892), .ZN(n1660) );
  aoi22d1 U2385 ( .A1(\RegFilePlugin_regFile[25][18] ), .A2(n1926), .B1(
        \RegFilePlugin_regFile[15][18] ), .B2(n1994), .ZN(n1659) );
  aoi22d1 U2386 ( .A1(\RegFilePlugin_regFile[20][18] ), .A2(n1387), .B1(
        \RegFilePlugin_regFile[19][18] ), .B2(n2024), .ZN(n1658) );
  aoi22d1 U2387 ( .A1(\RegFilePlugin_regFile[5][18] ), .A2(n1982), .B1(
        \RegFilePlugin_regFile[13][18] ), .B2(n1932), .ZN(n1665) );
  aoi22d1 U2388 ( .A1(\RegFilePlugin_regFile[9][18] ), .A2(n1858), .B1(
        \RegFilePlugin_regFile[0][18] ), .B2(n2030), .ZN(n1664) );
  aoi22d1 U2389 ( .A1(\RegFilePlugin_regFile[27][18] ), .A2(n1718), .B1(
        \RegFilePlugin_regFile[10][18] ), .B2(n1416), .ZN(n1663) );
  aoi22d1 U2390 ( .A1(\RegFilePlugin_regFile[2][18] ), .A2(n2032), .B1(
        \RegFilePlugin_regFile[30][18] ), .B2(n1987), .ZN(n1662) );
  or04d0 U2391 ( .A1(n1669), .A2(n1668), .A3(n1667), .A4(n1666), .Z(N869) );
  aoi22d1 U2392 ( .A1(\RegFilePlugin_regFile[10][16] ), .A2(n1416), .B1(
        \RegFilePlugin_regFile[24][16] ), .B2(n1735), .ZN(n1675) );
  aoi22d1 U2393 ( .A1(\RegFilePlugin_regFile[8][16] ), .A2(n1670), .B1(
        \RegFilePlugin_regFile[18][16] ), .B2(n1937), .ZN(n1674) );
  aoi22d1 U2394 ( .A1(\RegFilePlugin_regFile[16][16] ), .A2(n1671), .B1(
        \RegFilePlugin_regFile[1][16] ), .B2(n1692), .ZN(n1673) );
  aoi22d1 U2395 ( .A1(\RegFilePlugin_regFile[21][16] ), .A2(n1377), .B1(
        \RegFilePlugin_regFile[17][16] ), .B2(n1976), .ZN(n1672) );
  aoi22d1 U2396 ( .A1(\RegFilePlugin_regFile[25][16] ), .A2(n1607), .B1(
        \RegFilePlugin_regFile[11][16] ), .B2(n2013), .ZN(n1679) );
  aoi22d1 U2397 ( .A1(\RegFilePlugin_regFile[22][16] ), .A2(n2014), .B1(
        \RegFilePlugin_regFile[9][16] ), .B2(n1858), .ZN(n1678) );
  aoi22d1 U2398 ( .A1(\RegFilePlugin_regFile[4][16] ), .A2(n2004), .B1(
        \RegFilePlugin_regFile[15][16] ), .B2(n1994), .ZN(n1677) );
  aoi22d1 U2399 ( .A1(\RegFilePlugin_regFile[12][16] ), .A2(n2031), .B1(
        \RegFilePlugin_regFile[5][16] ), .B2(n1606), .ZN(n1676) );
  aoi22d1 U2400 ( .A1(\RegFilePlugin_regFile[13][16] ), .A2(n1932), .B1(
        \RegFilePlugin_regFile[0][16] ), .B2(n1585), .ZN(n1683) );
  aoi22d1 U2401 ( .A1(\RegFilePlugin_regFile[20][16] ), .A2(n1387), .B1(
        \RegFilePlugin_regFile[14][16] ), .B2(n1916), .ZN(n1682) );
  aoi22d1 U2402 ( .A1(\RegFilePlugin_regFile[7][16] ), .A2(n1543), .B1(
        \RegFilePlugin_regFile[6][16] ), .B2(n1943), .ZN(n1681) );
  aoi22d1 U2403 ( .A1(\RegFilePlugin_regFile[29][16] ), .A2(n1501), .B1(
        \RegFilePlugin_regFile[23][16] ), .B2(n2021), .ZN(n1680) );
  aoi22d1 U2404 ( .A1(\RegFilePlugin_regFile[3][16] ), .A2(n2022), .B1(
        \RegFilePlugin_regFile[26][16] ), .B2(n2015), .ZN(n1687) );
  aoi22d1 U2405 ( .A1(\RegFilePlugin_regFile[30][16] ), .A2(n1987), .B1(
        \RegFilePlugin_regFile[19][16] ), .B2(n1458), .ZN(n1686) );
  aoi22d1 U2406 ( .A1(\RegFilePlugin_regFile[27][16] ), .A2(n2033), .B1(
        \RegFilePlugin_regFile[2][16] ), .B2(n1628), .ZN(n1685) );
  aoi22d1 U2407 ( .A1(\RegFilePlugin_regFile[31][16] ), .A2(n1417), .B1(
        \RegFilePlugin_regFile[28][16] ), .B2(n1892), .ZN(n1684) );
  or04d0 U2408 ( .A1(n1691), .A2(n1690), .A3(n1689), .A4(n1688), .Z(N871) );
  aoi22d1 U2409 ( .A1(\RegFilePlugin_regFile[1][7] ), .A2(n1692), .B1(
        \RegFilePlugin_regFile[29][7] ), .B2(n1974), .ZN(n1696) );
  aoi22d1 U2410 ( .A1(\RegFilePlugin_regFile[31][7] ), .A2(n1417), .B1(
        \RegFilePlugin_regFile[12][7] ), .B2(n1981), .ZN(n1695) );
  aoi22d1 U2411 ( .A1(\RegFilePlugin_regFile[10][7] ), .A2(n1993), .B1(
        \RegFilePlugin_regFile[2][7] ), .B2(n1628), .ZN(n1694) );
  aoi22d1 U2412 ( .A1(\RegFilePlugin_regFile[6][7] ), .A2(n1522), .B1(
        \RegFilePlugin_regFile[30][7] ), .B2(n1987), .ZN(n1693) );
  aoi22d1 U2413 ( .A1(\RegFilePlugin_regFile[5][7] ), .A2(n1982), .B1(
        \RegFilePlugin_regFile[17][7] ), .B2(n1976), .ZN(n1701) );
  aoi22d1 U2414 ( .A1(\RegFilePlugin_regFile[15][7] ), .A2(n1697), .B1(
        \RegFilePlugin_regFile[0][7] ), .B2(n2030), .ZN(n1700) );
  aoi22d1 U2415 ( .A1(\RegFilePlugin_regFile[28][7] ), .A2(n1903), .B1(
        \RegFilePlugin_regFile[3][7] ), .B2(n2022), .ZN(n1699) );
  aoi22d1 U2416 ( .A1(\RegFilePlugin_regFile[19][7] ), .A2(n2024), .B1(
        \RegFilePlugin_regFile[4][7] ), .B2(n2004), .ZN(n1698) );
  aoi22d1 U2417 ( .A1(\RegFilePlugin_regFile[25][7] ), .A2(n1607), .B1(
        \RegFilePlugin_regFile[27][7] ), .B2(n1718), .ZN(n1705) );
  aoi22d1 U2418 ( .A1(\RegFilePlugin_regFile[24][7] ), .A2(n1735), .B1(
        \RegFilePlugin_regFile[13][7] ), .B2(n1932), .ZN(n1704) );
  aoi22d1 U2419 ( .A1(\RegFilePlugin_regFile[18][7] ), .A2(n1937), .B1(
        \RegFilePlugin_regFile[20][7] ), .B2(n2006), .ZN(n1703) );
  aoi22d1 U2420 ( .A1(\RegFilePlugin_regFile[26][7] ), .A2(n2015), .B1(
        \RegFilePlugin_regFile[21][7] ), .B2(n1931), .ZN(n1702) );
  aoi22d1 U2421 ( .A1(\RegFilePlugin_regFile[22][7] ), .A2(n2014), .B1(
        \RegFilePlugin_regFile[7][7] ), .B2(n1925), .ZN(n1709) );
  aoi22d1 U2422 ( .A1(\RegFilePlugin_regFile[8][7] ), .A2(n1902), .B1(
        \RegFilePlugin_regFile[9][7] ), .B2(n2011), .ZN(n1708) );
  aoi22d1 U2423 ( .A1(\RegFilePlugin_regFile[14][7] ), .A2(n2003), .B1(
        \RegFilePlugin_regFile[11][7] ), .B2(n2013), .ZN(n1707) );
  aoi22d1 U2424 ( .A1(\RegFilePlugin_regFile[23][7] ), .A2(n1544), .B1(
        \RegFilePlugin_regFile[16][7] ), .B2(n1975), .ZN(n1706) );
  or04d0 U2425 ( .A1(n1713), .A2(n1712), .A3(n1711), .A4(n1710), .Z(N880) );
  aoi22d1 U2426 ( .A1(\RegFilePlugin_regFile[10][10] ), .A2(n1993), .B1(
        \RegFilePlugin_regFile[21][10] ), .B2(n1377), .ZN(n1717) );
  aoi22d1 U2427 ( .A1(\RegFilePlugin_regFile[16][10] ), .A2(n1975), .B1(
        \RegFilePlugin_regFile[30][10] ), .B2(n1837), .ZN(n1716) );
  aoi22d1 U2428 ( .A1(\RegFilePlugin_regFile[31][10] ), .A2(n1417), .B1(
        \RegFilePlugin_regFile[24][10] ), .B2(n1735), .ZN(n1715) );
  aoi22d1 U2429 ( .A1(\RegFilePlugin_regFile[26][10] ), .A2(n2015), .B1(
        \RegFilePlugin_regFile[20][10] ), .B2(n2006), .ZN(n1714) );
  aoi22d1 U2430 ( .A1(\RegFilePlugin_regFile[3][10] ), .A2(n2022), .B1(
        \RegFilePlugin_regFile[29][10] ), .B2(n1501), .ZN(n1722) );
  aoi22d1 U2431 ( .A1(\RegFilePlugin_regFile[27][10] ), .A2(n1718), .B1(
        \RegFilePlugin_regFile[4][10] ), .B2(n2004), .ZN(n1721) );
  aoi22d1 U2432 ( .A1(\RegFilePlugin_regFile[9][10] ), .A2(n2011), .B1(
        \RegFilePlugin_regFile[23][10] ), .B2(n2021), .ZN(n1720) );
  aoi22d1 U2433 ( .A1(\RegFilePlugin_regFile[11][10] ), .A2(n2013), .B1(
        \RegFilePlugin_regFile[5][10] ), .B2(n1982), .ZN(n1719) );
  aoi22d1 U2434 ( .A1(\RegFilePlugin_regFile[12][10] ), .A2(n2031), .B1(
        \RegFilePlugin_regFile[25][10] ), .B2(n1926), .ZN(n1726) );
  aoi22d1 U2435 ( .A1(\RegFilePlugin_regFile[7][10] ), .A2(n1925), .B1(
        \RegFilePlugin_regFile[14][10] ), .B2(n2003), .ZN(n1725) );
  aoi22d1 U2436 ( .A1(\RegFilePlugin_regFile[8][10] ), .A2(n1670), .B1(
        \RegFilePlugin_regFile[2][10] ), .B2(n2032), .ZN(n1724) );
  aoi22d1 U2437 ( .A1(\RegFilePlugin_regFile[19][10] ), .A2(n2024), .B1(
        \RegFilePlugin_regFile[17][10] ), .B2(n1976), .ZN(n1723) );
  aoi22d1 U2438 ( .A1(\RegFilePlugin_regFile[22][10] ), .A2(n2014), .B1(
        \RegFilePlugin_regFile[1][10] ), .B2(n1692), .ZN(n1730) );
  aoi22d1 U2439 ( .A1(\RegFilePlugin_regFile[15][10] ), .A2(n2023), .B1(
        \RegFilePlugin_regFile[18][10] ), .B2(n1937), .ZN(n1729) );
  aoi22d1 U2440 ( .A1(\RegFilePlugin_regFile[0][10] ), .A2(n2030), .B1(
        \RegFilePlugin_regFile[6][10] ), .B2(n1943), .ZN(n1728) );
  aoi22d1 U2441 ( .A1(\RegFilePlugin_regFile[28][10] ), .A2(n1892), .B1(
        \RegFilePlugin_regFile[13][10] ), .B2(n2025), .ZN(n1727) );
  or04d0 U2442 ( .A1(n1734), .A2(n1733), .A3(n1732), .A4(n1731), .Z(N877) );
  aoi22d1 U2443 ( .A1(\RegFilePlugin_regFile[30][14] ), .A2(n1987), .B1(
        \RegFilePlugin_regFile[6][14] ), .B2(n1943), .ZN(n1739) );
  aoi22d1 U2444 ( .A1(\RegFilePlugin_regFile[19][14] ), .A2(n1458), .B1(
        \RegFilePlugin_regFile[24][14] ), .B2(n1735), .ZN(n1738) );
  aoi22d1 U2445 ( .A1(\RegFilePlugin_regFile[11][14] ), .A2(n1901), .B1(
        \RegFilePlugin_regFile[2][14] ), .B2(n1628), .ZN(n1737) );
  aoi22d1 U2446 ( .A1(\RegFilePlugin_regFile[12][14] ), .A2(n2031), .B1(
        \RegFilePlugin_regFile[5][14] ), .B2(n1606), .ZN(n1736) );
  aoi22d1 U2447 ( .A1(\RegFilePlugin_regFile[16][14] ), .A2(n1671), .B1(
        \RegFilePlugin_regFile[20][14] ), .B2(n2006), .ZN(n1743) );
  aoi22d1 U2448 ( .A1(\RegFilePlugin_regFile[10][14] ), .A2(n1416), .B1(
        \RegFilePlugin_regFile[26][14] ), .B2(n2015), .ZN(n1742) );
  aoi22d1 U2449 ( .A1(\RegFilePlugin_regFile[9][14] ), .A2(n1858), .B1(
        \RegFilePlugin_regFile[29][14] ), .B2(n1974), .ZN(n1741) );
  aoi22d1 U2450 ( .A1(\RegFilePlugin_regFile[0][14] ), .A2(n1585), .B1(
        \RegFilePlugin_regFile[22][14] ), .B2(n1988), .ZN(n1740) );
  aoi22d1 U2451 ( .A1(\RegFilePlugin_regFile[27][14] ), .A2(n2033), .B1(
        \RegFilePlugin_regFile[23][14] ), .B2(n2021), .ZN(n1747) );
  aoi22d1 U2452 ( .A1(\RegFilePlugin_regFile[17][14] ), .A2(n1976), .B1(
        \RegFilePlugin_regFile[28][14] ), .B2(n1892), .ZN(n1746) );
  aoi22d1 U2453 ( .A1(\RegFilePlugin_regFile[15][14] ), .A2(n1994), .B1(
        \RegFilePlugin_regFile[25][14] ), .B2(n1926), .ZN(n1745) );
  aoi22d1 U2454 ( .A1(\RegFilePlugin_regFile[3][14] ), .A2(n1816), .B1(
        \RegFilePlugin_regFile[21][14] ), .B2(n1377), .ZN(n1744) );
  aoi22d1 U2455 ( .A1(\RegFilePlugin_regFile[8][14] ), .A2(n1902), .B1(
        \RegFilePlugin_regFile[1][14] ), .B2(n1692), .ZN(n1751) );
  aoi22d1 U2456 ( .A1(\RegFilePlugin_regFile[13][14] ), .A2(n1932), .B1(
        \RegFilePlugin_regFile[14][14] ), .B2(n1916), .ZN(n1750) );
  aoi22d1 U2457 ( .A1(\RegFilePlugin_regFile[18][14] ), .A2(n1952), .B1(
        \RegFilePlugin_regFile[4][14] ), .B2(n2004), .ZN(n1749) );
  aoi22d1 U2458 ( .A1(\RegFilePlugin_regFile[7][14] ), .A2(n1543), .B1(
        \RegFilePlugin_regFile[31][14] ), .B2(n1942), .ZN(n1748) );
  or04d0 U2459 ( .A1(n1755), .A2(n1754), .A3(n1753), .A4(n1752), .Z(N873) );
  aoi22d1 U2460 ( .A1(\RegFilePlugin_regFile[30][22] ), .A2(n1837), .B1(
        \RegFilePlugin_regFile[26][22] ), .B2(n2015), .ZN(n1759) );
  aoi22d1 U2461 ( .A1(\RegFilePlugin_regFile[6][22] ), .A2(n1943), .B1(
        \RegFilePlugin_regFile[15][22] ), .B2(n2023), .ZN(n1758) );
  aoi22d1 U2462 ( .A1(\RegFilePlugin_regFile[13][22] ), .A2(n1932), .B1(
        \RegFilePlugin_regFile[27][22] ), .B2(n1718), .ZN(n1757) );
  aoi22d1 U2463 ( .A1(\RegFilePlugin_regFile[3][22] ), .A2(n1816), .B1(
        \RegFilePlugin_regFile[10][22] ), .B2(n1416), .ZN(n1756) );
  aoi22d1 U2464 ( .A1(\RegFilePlugin_regFile[19][22] ), .A2(n2024), .B1(
        \RegFilePlugin_regFile[14][22] ), .B2(n1916), .ZN(n1763) );
  aoi22d1 U2465 ( .A1(\RegFilePlugin_regFile[7][22] ), .A2(n1543), .B1(
        \RegFilePlugin_regFile[23][22] ), .B2(n2021), .ZN(n1762) );
  aoi22d1 U2466 ( .A1(\RegFilePlugin_regFile[28][22] ), .A2(n1892), .B1(
        \RegFilePlugin_regFile[22][22] ), .B2(n2014), .ZN(n1761) );
  aoi22d1 U2467 ( .A1(\RegFilePlugin_regFile[1][22] ), .A2(n2012), .B1(
        \RegFilePlugin_regFile[12][22] ), .B2(n1981), .ZN(n1760) );
  aoi22d1 U2468 ( .A1(\RegFilePlugin_regFile[31][22] ), .A2(n1942), .B1(
        \RegFilePlugin_regFile[29][22] ), .B2(n1974), .ZN(n1767) );
  aoi22d1 U2469 ( .A1(\RegFilePlugin_regFile[4][22] ), .A2(n1879), .B1(
        \RegFilePlugin_regFile[16][22] ), .B2(n1671), .ZN(n1766) );
  aoi22d1 U2470 ( .A1(\RegFilePlugin_regFile[11][22] ), .A2(n1901), .B1(
        \RegFilePlugin_regFile[18][22] ), .B2(n1937), .ZN(n1765) );
  aoi22d1 U2471 ( .A1(\RegFilePlugin_regFile[25][22] ), .A2(n1607), .B1(
        \RegFilePlugin_regFile[5][22] ), .B2(n1982), .ZN(n1764) );
  aoi22d1 U2472 ( .A1(\RegFilePlugin_regFile[21][22] ), .A2(n1377), .B1(
        \RegFilePlugin_regFile[0][22] ), .B2(n2030), .ZN(n1771) );
  aoi22d1 U2473 ( .A1(\RegFilePlugin_regFile[2][22] ), .A2(n2032), .B1(
        \RegFilePlugin_regFile[17][22] ), .B2(n1953), .ZN(n1770) );
  aoi22d1 U2474 ( .A1(\RegFilePlugin_regFile[8][22] ), .A2(n1902), .B1(
        \RegFilePlugin_regFile[20][22] ), .B2(n2006), .ZN(n1769) );
  aoi22d1 U2475 ( .A1(\RegFilePlugin_regFile[24][22] ), .A2(n2020), .B1(
        \RegFilePlugin_regFile[9][22] ), .B2(n1858), .ZN(n1768) );
  or04d0 U2476 ( .A1(n1775), .A2(n1774), .A3(n1773), .A4(n1772), .Z(N865) );
  aoi22d1 U2477 ( .A1(\RegFilePlugin_regFile[6][31] ), .A2(n1943), .B1(
        \RegFilePlugin_regFile[24][31] ), .B2(n2020), .ZN(n1779) );
  aoi22d1 U2478 ( .A1(\RegFilePlugin_regFile[25][31] ), .A2(n1926), .B1(
        \RegFilePlugin_regFile[29][31] ), .B2(n1501), .ZN(n1778) );
  aoi22d1 U2479 ( .A1(\RegFilePlugin_regFile[17][31] ), .A2(n1976), .B1(
        \RegFilePlugin_regFile[4][31] ), .B2(n1879), .ZN(n1777) );
  aoi22d1 U2480 ( .A1(\RegFilePlugin_regFile[22][31] ), .A2(n1988), .B1(
        \RegFilePlugin_regFile[5][31] ), .B2(n1606), .ZN(n1776) );
  aoi22d1 U2481 ( .A1(\RegFilePlugin_regFile[8][31] ), .A2(n1902), .B1(
        \RegFilePlugin_regFile[9][31] ), .B2(n1858), .ZN(n1783) );
  aoi22d1 U2482 ( .A1(\RegFilePlugin_regFile[19][31] ), .A2(n1458), .B1(
        \RegFilePlugin_regFile[16][31] ), .B2(n1975), .ZN(n1782) );
  aoi22d1 U2483 ( .A1(\RegFilePlugin_regFile[21][31] ), .A2(n1931), .B1(
        \RegFilePlugin_regFile[31][31] ), .B2(n1417), .ZN(n1781) );
  aoi22d1 U2484 ( .A1(\RegFilePlugin_regFile[26][31] ), .A2(n1649), .B1(
        \RegFilePlugin_regFile[14][31] ), .B2(n2003), .ZN(n1780) );
  aoi22d1 U2485 ( .A1(\RegFilePlugin_regFile[20][31] ), .A2(n2006), .B1(
        \RegFilePlugin_regFile[12][31] ), .B2(n1981), .ZN(n1787) );
  aoi22d1 U2486 ( .A1(\RegFilePlugin_regFile[3][31] ), .A2(n1816), .B1(
        \RegFilePlugin_regFile[28][31] ), .B2(n1903), .ZN(n1786) );
  aoi22d1 U2487 ( .A1(\RegFilePlugin_regFile[30][31] ), .A2(n1987), .B1(
        \RegFilePlugin_regFile[0][31] ), .B2(n1585), .ZN(n1785) );
  aoi22d1 U2488 ( .A1(\RegFilePlugin_regFile[1][31] ), .A2(n2012), .B1(
        \RegFilePlugin_regFile[23][31] ), .B2(n1544), .ZN(n1784) );
  aoi22d1 U2489 ( .A1(\RegFilePlugin_regFile[2][31] ), .A2(n1628), .B1(
        \RegFilePlugin_regFile[7][31] ), .B2(n1543), .ZN(n1791) );
  aoi22d1 U2490 ( .A1(\RegFilePlugin_regFile[10][31] ), .A2(n1993), .B1(
        \RegFilePlugin_regFile[15][31] ), .B2(n2023), .ZN(n1790) );
  aoi22d1 U2491 ( .A1(\RegFilePlugin_regFile[18][31] ), .A2(n1952), .B1(
        \RegFilePlugin_regFile[11][31] ), .B2(n1901), .ZN(n1789) );
  aoi22d1 U2492 ( .A1(\RegFilePlugin_regFile[13][31] ), .A2(n2025), .B1(
        \RegFilePlugin_regFile[27][31] ), .B2(n2033), .ZN(n1788) );
  or04d0 U2493 ( .A1(n1795), .A2(n1794), .A3(n1793), .A4(n1792), .Z(N856) );
  aoi22d1 U2494 ( .A1(\RegFilePlugin_regFile[8][13] ), .A2(n1670), .B1(
        \RegFilePlugin_regFile[4][13] ), .B2(n2004), .ZN(n1799) );
  aoi22d1 U2495 ( .A1(\RegFilePlugin_regFile[21][13] ), .A2(n1931), .B1(
        \RegFilePlugin_regFile[17][13] ), .B2(n1953), .ZN(n1798) );
  aoi22d1 U2496 ( .A1(\RegFilePlugin_regFile[29][13] ), .A2(n1974), .B1(
        \RegFilePlugin_regFile[3][13] ), .B2(n1816), .ZN(n1797) );
  aoi22d1 U2497 ( .A1(\RegFilePlugin_regFile[2][13] ), .A2(n2032), .B1(
        \RegFilePlugin_regFile[24][13] ), .B2(n1735), .ZN(n1796) );
  aoi22d1 U2498 ( .A1(\RegFilePlugin_regFile[6][13] ), .A2(n1943), .B1(
        \RegFilePlugin_regFile[5][13] ), .B2(n1606), .ZN(n1803) );
  aoi22d1 U2499 ( .A1(\RegFilePlugin_regFile[15][13] ), .A2(n1994), .B1(
        \RegFilePlugin_regFile[19][13] ), .B2(n1458), .ZN(n1802) );
  aoi22d1 U2500 ( .A1(\RegFilePlugin_regFile[31][13] ), .A2(n1417), .B1(
        \RegFilePlugin_regFile[0][13] ), .B2(n1585), .ZN(n1801) );
  aoi22d1 U2501 ( .A1(\RegFilePlugin_regFile[16][13] ), .A2(n1975), .B1(
        \RegFilePlugin_regFile[30][13] ), .B2(n1837), .ZN(n1800) );
  aoi22d1 U2502 ( .A1(\RegFilePlugin_regFile[12][13] ), .A2(n2031), .B1(
        \RegFilePlugin_regFile[28][13] ), .B2(n1892), .ZN(n1807) );
  aoi22d1 U2503 ( .A1(\RegFilePlugin_regFile[27][13] ), .A2(n1718), .B1(
        \RegFilePlugin_regFile[11][13] ), .B2(n2013), .ZN(n1806) );
  aoi22d1 U2504 ( .A1(\RegFilePlugin_regFile[9][13] ), .A2(n2011), .B1(
        \RegFilePlugin_regFile[23][13] ), .B2(n1544), .ZN(n1805) );
  aoi22d1 U2505 ( .A1(\RegFilePlugin_regFile[22][13] ), .A2(n1988), .B1(
        \RegFilePlugin_regFile[18][13] ), .B2(n1937), .ZN(n1804) );
  aoi22d1 U2506 ( .A1(\RegFilePlugin_regFile[20][13] ), .A2(n1387), .B1(
        \RegFilePlugin_regFile[26][13] ), .B2(n2015), .ZN(n1811) );
  aoi22d1 U2507 ( .A1(\RegFilePlugin_regFile[25][13] ), .A2(n1607), .B1(
        \RegFilePlugin_regFile[10][13] ), .B2(n1416), .ZN(n1810) );
  aoi22d1 U2508 ( .A1(\RegFilePlugin_regFile[13][13] ), .A2(n2025), .B1(
        \RegFilePlugin_regFile[1][13] ), .B2(n1692), .ZN(n1809) );
  aoi22d1 U2509 ( .A1(\RegFilePlugin_regFile[14][13] ), .A2(n2003), .B1(
        \RegFilePlugin_regFile[7][13] ), .B2(n1925), .ZN(n1808) );
  or04d0 U2510 ( .A1(n1815), .A2(n1814), .A3(n1813), .A4(n1812), .Z(N874) );
  aoi22d1 U2511 ( .A1(\RegFilePlugin_regFile[5][1] ), .A2(n1606), .B1(
        \RegFilePlugin_regFile[0][1] ), .B2(n1585), .ZN(n1820) );
  aoi22d1 U2512 ( .A1(\RegFilePlugin_regFile[25][1] ), .A2(n1926), .B1(
        \RegFilePlugin_regFile[1][1] ), .B2(n2012), .ZN(n1819) );
  aoi22d1 U2513 ( .A1(\RegFilePlugin_regFile[31][1] ), .A2(n1417), .B1(
        \RegFilePlugin_regFile[9][1] ), .B2(n2011), .ZN(n1818) );
  aoi22d1 U2514 ( .A1(\RegFilePlugin_regFile[3][1] ), .A2(n1816), .B1(
        \RegFilePlugin_regFile[20][1] ), .B2(n1387), .ZN(n1817) );
  aoi22d1 U2515 ( .A1(\RegFilePlugin_regFile[26][1] ), .A2(n1649), .B1(
        \RegFilePlugin_regFile[15][1] ), .B2(n1994), .ZN(n1824) );
  aoi22d1 U2516 ( .A1(\RegFilePlugin_regFile[19][1] ), .A2(n2024), .B1(
        \RegFilePlugin_regFile[29][1] ), .B2(n1501), .ZN(n1823) );
  aoi22d1 U2517 ( .A1(\RegFilePlugin_regFile[28][1] ), .A2(n1903), .B1(
        \RegFilePlugin_regFile[22][1] ), .B2(n1988), .ZN(n1822) );
  aoi22d1 U2518 ( .A1(\RegFilePlugin_regFile[27][1] ), .A2(n2033), .B1(
        \RegFilePlugin_regFile[10][1] ), .B2(n1993), .ZN(n1821) );
  aoi22d1 U2519 ( .A1(\RegFilePlugin_regFile[30][1] ), .A2(n1837), .B1(
        \RegFilePlugin_regFile[16][1] ), .B2(n1975), .ZN(n1828) );
  aoi22d1 U2520 ( .A1(\RegFilePlugin_regFile[17][1] ), .A2(n1976), .B1(
        \RegFilePlugin_regFile[4][1] ), .B2(n1879), .ZN(n1827) );
  aoi22d1 U2521 ( .A1(\RegFilePlugin_regFile[23][1] ), .A2(n2021), .B1(
        \RegFilePlugin_regFile[14][1] ), .B2(n1916), .ZN(n1826) );
  aoi22d1 U2522 ( .A1(\RegFilePlugin_regFile[12][1] ), .A2(n1981), .B1(
        \RegFilePlugin_regFile[7][1] ), .B2(n1543), .ZN(n1825) );
  aoi22d1 U2523 ( .A1(\RegFilePlugin_regFile[18][1] ), .A2(n1937), .B1(
        \RegFilePlugin_regFile[11][1] ), .B2(n2013), .ZN(n1832) );
  aoi22d1 U2524 ( .A1(\RegFilePlugin_regFile[2][1] ), .A2(n2032), .B1(
        \RegFilePlugin_regFile[21][1] ), .B2(n1377), .ZN(n1831) );
  aoi22d1 U2525 ( .A1(\RegFilePlugin_regFile[6][1] ), .A2(n1522), .B1(
        \RegFilePlugin_regFile[24][1] ), .B2(n1735), .ZN(n1830) );
  aoi22d1 U2526 ( .A1(\RegFilePlugin_regFile[13][1] ), .A2(n2025), .B1(
        \RegFilePlugin_regFile[8][1] ), .B2(n1670), .ZN(n1829) );
  or04d0 U2527 ( .A1(n1836), .A2(n1835), .A3(n1834), .A4(n1833), .Z(N886) );
  aoi22d1 U2528 ( .A1(\RegFilePlugin_regFile[30][8] ), .A2(n1837), .B1(
        \RegFilePlugin_regFile[8][8] ), .B2(n1670), .ZN(n1841) );
  aoi22d1 U2529 ( .A1(\RegFilePlugin_regFile[27][8] ), .A2(n1718), .B1(
        \RegFilePlugin_regFile[23][8] ), .B2(n1544), .ZN(n1840) );
  aoi22d1 U2530 ( .A1(\RegFilePlugin_regFile[6][8] ), .A2(n1522), .B1(
        \RegFilePlugin_regFile[22][8] ), .B2(n1988), .ZN(n1839) );
  aoi22d1 U2531 ( .A1(\RegFilePlugin_regFile[17][8] ), .A2(n1976), .B1(
        \RegFilePlugin_regFile[15][8] ), .B2(n1994), .ZN(n1838) );
  aoi22d1 U2532 ( .A1(\RegFilePlugin_regFile[13][8] ), .A2(n1932), .B1(
        \RegFilePlugin_regFile[3][8] ), .B2(n2022), .ZN(n1845) );
  aoi22d1 U2533 ( .A1(\RegFilePlugin_regFile[14][8] ), .A2(n2003), .B1(
        \RegFilePlugin_regFile[12][8] ), .B2(n1981), .ZN(n1844) );
  aoi22d1 U2534 ( .A1(\RegFilePlugin_regFile[7][8] ), .A2(n1925), .B1(
        \RegFilePlugin_regFile[11][8] ), .B2(n1901), .ZN(n1843) );
  aoi22d1 U2535 ( .A1(\RegFilePlugin_regFile[25][8] ), .A2(n1607), .B1(
        \RegFilePlugin_regFile[0][8] ), .B2(n1585), .ZN(n1842) );
  aoi22d1 U2536 ( .A1(\RegFilePlugin_regFile[19][8] ), .A2(n1458), .B1(
        \RegFilePlugin_regFile[5][8] ), .B2(n1982), .ZN(n1849) );
  aoi22d1 U2537 ( .A1(\RegFilePlugin_regFile[28][8] ), .A2(n1903), .B1(
        \RegFilePlugin_regFile[31][8] ), .B2(n1942), .ZN(n1848) );
  aoi22d1 U2538 ( .A1(\RegFilePlugin_regFile[4][8] ), .A2(n1879), .B1(
        \RegFilePlugin_regFile[10][8] ), .B2(n1993), .ZN(n1847) );
  aoi22d1 U2539 ( .A1(\RegFilePlugin_regFile[16][8] ), .A2(n1975), .B1(
        \RegFilePlugin_regFile[29][8] ), .B2(n1974), .ZN(n1846) );
  aoi22d1 U2540 ( .A1(\RegFilePlugin_regFile[21][8] ), .A2(n1931), .B1(
        \RegFilePlugin_regFile[2][8] ), .B2(n1628), .ZN(n1853) );
  aoi22d1 U2541 ( .A1(\RegFilePlugin_regFile[1][8] ), .A2(n2012), .B1(
        \RegFilePlugin_regFile[9][8] ), .B2(n1858), .ZN(n1852) );
  aoi22d1 U2542 ( .A1(\RegFilePlugin_regFile[18][8] ), .A2(n1952), .B1(
        \RegFilePlugin_regFile[24][8] ), .B2(n2020), .ZN(n1851) );
  aoi22d1 U2543 ( .A1(\RegFilePlugin_regFile[26][8] ), .A2(n1649), .B1(
        \RegFilePlugin_regFile[20][8] ), .B2(n1387), .ZN(n1850) );
  or04d0 U2544 ( .A1(n1857), .A2(n1856), .A3(n1855), .A4(n1854), .Z(N879) );
  aoi22d1 U2545 ( .A1(\RegFilePlugin_regFile[9][17] ), .A2(n1858), .B1(
        \RegFilePlugin_regFile[3][17] ), .B2(n2022), .ZN(n1862) );
  aoi22d1 U2546 ( .A1(\RegFilePlugin_regFile[12][17] ), .A2(n2031), .B1(
        \RegFilePlugin_regFile[18][17] ), .B2(n1952), .ZN(n1861) );
  aoi22d1 U2547 ( .A1(\RegFilePlugin_regFile[4][17] ), .A2(n1879), .B1(
        \RegFilePlugin_regFile[5][17] ), .B2(n1606), .ZN(n1860) );
  aoi22d1 U2548 ( .A1(\RegFilePlugin_regFile[30][17] ), .A2(n1987), .B1(
        \RegFilePlugin_regFile[24][17] ), .B2(n2020), .ZN(n1859) );
  aoi22d1 U2549 ( .A1(\RegFilePlugin_regFile[6][17] ), .A2(n1522), .B1(
        \RegFilePlugin_regFile[31][17] ), .B2(n1942), .ZN(n1866) );
  aoi22d1 U2550 ( .A1(\RegFilePlugin_regFile[23][17] ), .A2(n2021), .B1(
        \RegFilePlugin_regFile[8][17] ), .B2(n1670), .ZN(n1865) );
  aoi22d1 U2551 ( .A1(\RegFilePlugin_regFile[2][17] ), .A2(n2032), .B1(
        \RegFilePlugin_regFile[22][17] ), .B2(n1988), .ZN(n1864) );
  aoi22d1 U2552 ( .A1(\RegFilePlugin_regFile[25][17] ), .A2(n1926), .B1(
        \RegFilePlugin_regFile[14][17] ), .B2(n1916), .ZN(n1863) );
  aoi22d1 U2553 ( .A1(\RegFilePlugin_regFile[27][17] ), .A2(n2033), .B1(
        \RegFilePlugin_regFile[26][17] ), .B2(n2015), .ZN(n1870) );
  aoi22d1 U2554 ( .A1(\RegFilePlugin_regFile[17][17] ), .A2(n1976), .B1(
        \RegFilePlugin_regFile[10][17] ), .B2(n1416), .ZN(n1869) );
  aoi22d1 U2555 ( .A1(\RegFilePlugin_regFile[20][17] ), .A2(n2006), .B1(
        \RegFilePlugin_regFile[1][17] ), .B2(n1692), .ZN(n1868) );
  aoi22d1 U2556 ( .A1(\RegFilePlugin_regFile[11][17] ), .A2(n1901), .B1(
        \RegFilePlugin_regFile[19][17] ), .B2(n1458), .ZN(n1867) );
  aoi22d1 U2557 ( .A1(\RegFilePlugin_regFile[7][17] ), .A2(n1925), .B1(
        \RegFilePlugin_regFile[29][17] ), .B2(n1974), .ZN(n1874) );
  aoi22d1 U2558 ( .A1(\RegFilePlugin_regFile[15][17] ), .A2(n1994), .B1(
        \RegFilePlugin_regFile[13][17] ), .B2(n1932), .ZN(n1873) );
  aoi22d1 U2559 ( .A1(\RegFilePlugin_regFile[16][17] ), .A2(n1671), .B1(
        \RegFilePlugin_regFile[28][17] ), .B2(n1892), .ZN(n1872) );
  aoi22d1 U2560 ( .A1(\RegFilePlugin_regFile[21][17] ), .A2(n1377), .B1(
        \RegFilePlugin_regFile[0][17] ), .B2(n2030), .ZN(n1871) );
  or04d0 U2561 ( .A1(n1878), .A2(n1877), .A3(n1876), .A4(n1875), .Z(N870) );
  aoi22d1 U2562 ( .A1(\RegFilePlugin_regFile[8][24] ), .A2(n1902), .B1(
        \RegFilePlugin_regFile[17][24] ), .B2(n1953), .ZN(n1883) );
  aoi22d1 U2563 ( .A1(\RegFilePlugin_regFile[4][24] ), .A2(n1879), .B1(
        \RegFilePlugin_regFile[13][24] ), .B2(n1932), .ZN(n1882) );
  aoi22d1 U2564 ( .A1(\RegFilePlugin_regFile[23][24] ), .A2(n1544), .B1(
        \RegFilePlugin_regFile[27][24] ), .B2(n1718), .ZN(n1881) );
  aoi22d1 U2565 ( .A1(\RegFilePlugin_regFile[3][24] ), .A2(n1816), .B1(
        \RegFilePlugin_regFile[16][24] ), .B2(n1671), .ZN(n1880) );
  aoi22d1 U2566 ( .A1(\RegFilePlugin_regFile[24][24] ), .A2(n2020), .B1(
        \RegFilePlugin_regFile[21][24] ), .B2(n1377), .ZN(n1887) );
  aoi22d1 U2567 ( .A1(\RegFilePlugin_regFile[12][24] ), .A2(n2031), .B1(
        \RegFilePlugin_regFile[30][24] ), .B2(n1837), .ZN(n1886) );
  aoi22d1 U2568 ( .A1(\RegFilePlugin_regFile[9][24] ), .A2(n2011), .B1(
        \RegFilePlugin_regFile[14][24] ), .B2(n1916), .ZN(n1885) );
  aoi22d1 U2569 ( .A1(\RegFilePlugin_regFile[15][24] ), .A2(n1994), .B1(
        \RegFilePlugin_regFile[2][24] ), .B2(n1628), .ZN(n1884) );
  aoi22d1 U2570 ( .A1(\RegFilePlugin_regFile[20][24] ), .A2(n2006), .B1(
        \RegFilePlugin_regFile[1][24] ), .B2(n1692), .ZN(n1891) );
  aoi22d1 U2571 ( .A1(\RegFilePlugin_regFile[6][24] ), .A2(n1943), .B1(
        \RegFilePlugin_regFile[29][24] ), .B2(n1501), .ZN(n1890) );
  aoi22d1 U2572 ( .A1(\RegFilePlugin_regFile[11][24] ), .A2(n1901), .B1(
        \RegFilePlugin_regFile[0][24] ), .B2(n1585), .ZN(n1889) );
  aoi22d1 U2573 ( .A1(\RegFilePlugin_regFile[18][24] ), .A2(n1952), .B1(
        \RegFilePlugin_regFile[19][24] ), .B2(n1458), .ZN(n1888) );
  aoi22d1 U2574 ( .A1(\RegFilePlugin_regFile[7][24] ), .A2(n1543), .B1(
        \RegFilePlugin_regFile[22][24] ), .B2(n2014), .ZN(n1896) );
  aoi22d1 U2575 ( .A1(\RegFilePlugin_regFile[10][24] ), .A2(n1993), .B1(
        \RegFilePlugin_regFile[5][24] ), .B2(n1982), .ZN(n1895) );
  aoi22d1 U2576 ( .A1(\RegFilePlugin_regFile[25][24] ), .A2(n1926), .B1(
        \RegFilePlugin_regFile[31][24] ), .B2(n1942), .ZN(n1894) );
  aoi22d1 U2577 ( .A1(\RegFilePlugin_regFile[28][24] ), .A2(n1892), .B1(
        \RegFilePlugin_regFile[26][24] ), .B2(n2015), .ZN(n1893) );
  or04d0 U2578 ( .A1(n1900), .A2(n1899), .A3(n1898), .A4(n1897), .Z(N863) );
  aoi22d1 U2579 ( .A1(\RegFilePlugin_regFile[8][12] ), .A2(n1902), .B1(
        \RegFilePlugin_regFile[11][12] ), .B2(n1901), .ZN(n1907) );
  aoi22d1 U2580 ( .A1(\RegFilePlugin_regFile[10][12] ), .A2(n1416), .B1(
        \RegFilePlugin_regFile[1][12] ), .B2(n2012), .ZN(n1906) );
  aoi22d1 U2581 ( .A1(\RegFilePlugin_regFile[18][12] ), .A2(n1952), .B1(
        \RegFilePlugin_regFile[13][12] ), .B2(n1932), .ZN(n1905) );
  aoi22d1 U2582 ( .A1(\RegFilePlugin_regFile[24][12] ), .A2(n1735), .B1(
        \RegFilePlugin_regFile[28][12] ), .B2(n1903), .ZN(n1904) );
  aoi22d1 U2583 ( .A1(\RegFilePlugin_regFile[3][12] ), .A2(n2022), .B1(
        \RegFilePlugin_regFile[22][12] ), .B2(n1988), .ZN(n1911) );
  aoi22d1 U2584 ( .A1(\RegFilePlugin_regFile[25][12] ), .A2(n1607), .B1(
        \RegFilePlugin_regFile[26][12] ), .B2(n1649), .ZN(n1910) );
  aoi22d1 U2585 ( .A1(\RegFilePlugin_regFile[7][12] ), .A2(n1543), .B1(
        \RegFilePlugin_regFile[17][12] ), .B2(n1953), .ZN(n1909) );
  aoi22d1 U2586 ( .A1(\RegFilePlugin_regFile[29][12] ), .A2(n1974), .B1(
        \RegFilePlugin_regFile[31][12] ), .B2(n1417), .ZN(n1908) );
  aoi22d1 U2587 ( .A1(\RegFilePlugin_regFile[9][12] ), .A2(n2011), .B1(
        \RegFilePlugin_regFile[12][12] ), .B2(n1981), .ZN(n1915) );
  aoi22d1 U2588 ( .A1(\RegFilePlugin_regFile[21][12] ), .A2(n1931), .B1(
        \RegFilePlugin_regFile[30][12] ), .B2(n1987), .ZN(n1914) );
  aoi22d1 U2589 ( .A1(\RegFilePlugin_regFile[20][12] ), .A2(n1387), .B1(
        \RegFilePlugin_regFile[23][12] ), .B2(n1544), .ZN(n1913) );
  aoi22d1 U2590 ( .A1(\RegFilePlugin_regFile[19][12] ), .A2(n2024), .B1(
        \RegFilePlugin_regFile[16][12] ), .B2(n1671), .ZN(n1912) );
  aoi22d1 U2591 ( .A1(\RegFilePlugin_regFile[5][12] ), .A2(n1982), .B1(
        \RegFilePlugin_regFile[14][12] ), .B2(n1916), .ZN(n1920) );
  aoi22d1 U2592 ( .A1(\RegFilePlugin_regFile[6][12] ), .A2(n1943), .B1(
        \RegFilePlugin_regFile[0][12] ), .B2(n1585), .ZN(n1919) );
  aoi22d1 U2593 ( .A1(\RegFilePlugin_regFile[4][12] ), .A2(n1879), .B1(
        \RegFilePlugin_regFile[15][12] ), .B2(n1994), .ZN(n1918) );
  aoi22d1 U2594 ( .A1(\RegFilePlugin_regFile[27][12] ), .A2(n2033), .B1(
        \RegFilePlugin_regFile[2][12] ), .B2(n1628), .ZN(n1917) );
  or04d0 U2595 ( .A1(n1924), .A2(n1923), .A3(n1922), .A4(n1921), .Z(N875) );
  aoi22d1 U2596 ( .A1(\RegFilePlugin_regFile[8][11] ), .A2(n1670), .B1(
        \RegFilePlugin_regFile[0][11] ), .B2(n1585), .ZN(n1930) );
  aoi22d1 U2597 ( .A1(\RegFilePlugin_regFile[7][11] ), .A2(n1925), .B1(
        \RegFilePlugin_regFile[19][11] ), .B2(n1458), .ZN(n1929) );
  aoi22d1 U2598 ( .A1(\RegFilePlugin_regFile[12][11] ), .A2(n1981), .B1(
        \RegFilePlugin_regFile[25][11] ), .B2(n1926), .ZN(n1928) );
  aoi22d1 U2599 ( .A1(\RegFilePlugin_regFile[24][11] ), .A2(n1735), .B1(
        \RegFilePlugin_regFile[10][11] ), .B2(n1416), .ZN(n1927) );
  aoi22d1 U2600 ( .A1(\RegFilePlugin_regFile[4][11] ), .A2(n1879), .B1(
        \RegFilePlugin_regFile[20][11] ), .B2(n2006), .ZN(n1936) );
  aoi22d1 U2601 ( .A1(\RegFilePlugin_regFile[13][11] ), .A2(n1932), .B1(
        \RegFilePlugin_regFile[21][11] ), .B2(n1931), .ZN(n1935) );
  aoi22d1 U2602 ( .A1(\RegFilePlugin_regFile[28][11] ), .A2(n1903), .B1(
        \RegFilePlugin_regFile[22][11] ), .B2(n1988), .ZN(n1934) );
  aoi22d1 U2603 ( .A1(\RegFilePlugin_regFile[26][11] ), .A2(n1649), .B1(
        \RegFilePlugin_regFile[5][11] ), .B2(n1606), .ZN(n1933) );
  aoi22d1 U2604 ( .A1(\RegFilePlugin_regFile[3][11] ), .A2(n2022), .B1(
        \RegFilePlugin_regFile[18][11] ), .B2(n1937), .ZN(n1941) );
  aoi22d1 U2605 ( .A1(\RegFilePlugin_regFile[23][11] ), .A2(n1544), .B1(
        \RegFilePlugin_regFile[2][11] ), .B2(n1628), .ZN(n1940) );
  aoi22d1 U2606 ( .A1(\RegFilePlugin_regFile[17][11] ), .A2(n1976), .B1(
        \RegFilePlugin_regFile[29][11] ), .B2(n1974), .ZN(n1939) );
  aoi22d1 U2607 ( .A1(\RegFilePlugin_regFile[1][11] ), .A2(n2012), .B1(
        \RegFilePlugin_regFile[9][11] ), .B2(n1858), .ZN(n1938) );
  aoi22d1 U2608 ( .A1(\RegFilePlugin_regFile[15][11] ), .A2(n2023), .B1(
        \RegFilePlugin_regFile[11][11] ), .B2(n2013), .ZN(n1947) );
  aoi22d1 U2609 ( .A1(\RegFilePlugin_regFile[30][11] ), .A2(n1837), .B1(
        \RegFilePlugin_regFile[31][11] ), .B2(n1942), .ZN(n1946) );
  aoi22d1 U2610 ( .A1(\RegFilePlugin_regFile[14][11] ), .A2(n2003), .B1(
        \RegFilePlugin_regFile[6][11] ), .B2(n1943), .ZN(n1945) );
  aoi22d1 U2611 ( .A1(\RegFilePlugin_regFile[16][11] ), .A2(n1975), .B1(
        \RegFilePlugin_regFile[27][11] ), .B2(n1718), .ZN(n1944) );
  or04d0 U2612 ( .A1(n1951), .A2(n1950), .A3(n1949), .A4(n1948), .Z(N876) );
  aoi22d1 U2613 ( .A1(\RegFilePlugin_regFile[18][3] ), .A2(n1952), .B1(
        \RegFilePlugin_regFile[14][3] ), .B2(n2003), .ZN(n1957) );
  aoi22d1 U2614 ( .A1(\RegFilePlugin_regFile[3][3] ), .A2(n2022), .B1(
        \RegFilePlugin_regFile[29][3] ), .B2(n1974), .ZN(n1956) );
  aoi22d1 U2615 ( .A1(\RegFilePlugin_regFile[30][3] ), .A2(n1837), .B1(
        \RegFilePlugin_regFile[7][3] ), .B2(n1925), .ZN(n1955) );
  aoi22d1 U2616 ( .A1(\RegFilePlugin_regFile[17][3] ), .A2(n1953), .B1(
        \RegFilePlugin_regFile[20][3] ), .B2(n1387), .ZN(n1954) );
  aoi22d1 U2617 ( .A1(\RegFilePlugin_regFile[10][3] ), .A2(n1993), .B1(
        \RegFilePlugin_regFile[16][3] ), .B2(n1975), .ZN(n1961) );
  aoi22d1 U2618 ( .A1(\RegFilePlugin_regFile[23][3] ), .A2(n2021), .B1(
        \RegFilePlugin_regFile[9][3] ), .B2(n1858), .ZN(n1960) );
  aoi22d1 U2619 ( .A1(\RegFilePlugin_regFile[28][3] ), .A2(n1892), .B1(
        \RegFilePlugin_regFile[22][3] ), .B2(n2014), .ZN(n1959) );
  aoi22d1 U2620 ( .A1(\RegFilePlugin_regFile[25][3] ), .A2(n1926), .B1(
        \RegFilePlugin_regFile[11][3] ), .B2(n1901), .ZN(n1958) );
  aoi22d1 U2621 ( .A1(\RegFilePlugin_regFile[0][3] ), .A2(n2030), .B1(
        \RegFilePlugin_regFile[27][3] ), .B2(n2033), .ZN(n1965) );
  aoi22d1 U2622 ( .A1(\RegFilePlugin_regFile[5][3] ), .A2(n1982), .B1(
        \RegFilePlugin_regFile[6][3] ), .B2(n1522), .ZN(n1964) );
  aoi22d1 U2623 ( .A1(\RegFilePlugin_regFile[26][3] ), .A2(n2015), .B1(
        \RegFilePlugin_regFile[13][3] ), .B2(n2025), .ZN(n1963) );
  aoi22d1 U2624 ( .A1(\RegFilePlugin_regFile[31][3] ), .A2(n1417), .B1(
        \RegFilePlugin_regFile[12][3] ), .B2(n1981), .ZN(n1962) );
  aoi22d1 U2625 ( .A1(\RegFilePlugin_regFile[1][3] ), .A2(n2012), .B1(
        \RegFilePlugin_regFile[15][3] ), .B2(n2023), .ZN(n1969) );
  aoi22d1 U2626 ( .A1(\RegFilePlugin_regFile[8][3] ), .A2(n1902), .B1(
        \RegFilePlugin_regFile[4][3] ), .B2(n2004), .ZN(n1968) );
  aoi22d1 U2627 ( .A1(\RegFilePlugin_regFile[19][3] ), .A2(n1458), .B1(
        \RegFilePlugin_regFile[21][3] ), .B2(n1931), .ZN(n1967) );
  aoi22d1 U2628 ( .A1(\RegFilePlugin_regFile[24][3] ), .A2(n2020), .B1(
        \RegFilePlugin_regFile[2][3] ), .B2(n2032), .ZN(n1966) );
  or04d0 U2629 ( .A1(n1973), .A2(n1972), .A3(n1971), .A4(n1970), .Z(N884) );
  aoi22d1 U2630 ( .A1(\RegFilePlugin_regFile[16][2] ), .A2(n1975), .B1(
        \RegFilePlugin_regFile[29][2] ), .B2(n1974), .ZN(n1980) );
  aoi22d1 U2631 ( .A1(\RegFilePlugin_regFile[17][2] ), .A2(n1976), .B1(
        \RegFilePlugin_regFile[3][2] ), .B2(n2022), .ZN(n1979) );
  aoi22d1 U2632 ( .A1(\RegFilePlugin_regFile[8][2] ), .A2(n1670), .B1(
        \RegFilePlugin_regFile[21][2] ), .B2(n1377), .ZN(n1978) );
  aoi22d1 U2633 ( .A1(\RegFilePlugin_regFile[1][2] ), .A2(n1692), .B1(
        \RegFilePlugin_regFile[4][2] ), .B2(n1879), .ZN(n1977) );
  aoi22d1 U2634 ( .A1(\RegFilePlugin_regFile[13][2] ), .A2(n2025), .B1(
        \RegFilePlugin_regFile[12][2] ), .B2(n1981), .ZN(n1986) );
  aoi22d1 U2635 ( .A1(\RegFilePlugin_regFile[5][2] ), .A2(n1982), .B1(
        \RegFilePlugin_regFile[6][2] ), .B2(n1522), .ZN(n1985) );
  aoi22d1 U2636 ( .A1(\RegFilePlugin_regFile[19][2] ), .A2(n1458), .B1(
        \RegFilePlugin_regFile[31][2] ), .B2(n1417), .ZN(n1984) );
  aoi22d1 U2637 ( .A1(\RegFilePlugin_regFile[20][2] ), .A2(n2006), .B1(
        \RegFilePlugin_regFile[11][2] ), .B2(n1901), .ZN(n1983) );
  aoi22d1 U2638 ( .A1(\RegFilePlugin_regFile[22][2] ), .A2(n1988), .B1(
        \RegFilePlugin_regFile[30][2] ), .B2(n1987), .ZN(n1992) );
  aoi22d1 U2639 ( .A1(\RegFilePlugin_regFile[27][2] ), .A2(n2033), .B1(
        \RegFilePlugin_regFile[28][2] ), .B2(n1903), .ZN(n1991) );
  aoi22d1 U2640 ( .A1(\RegFilePlugin_regFile[0][2] ), .A2(n2030), .B1(
        \RegFilePlugin_regFile[9][2] ), .B2(n2011), .ZN(n1990) );
  aoi22d1 U2641 ( .A1(\RegFilePlugin_regFile[24][2] ), .A2(n1735), .B1(
        \RegFilePlugin_regFile[14][2] ), .B2(n2003), .ZN(n1989) );
  aoi22d1 U2642 ( .A1(\RegFilePlugin_regFile[2][2] ), .A2(n2032), .B1(
        \RegFilePlugin_regFile[7][2] ), .B2(n1543), .ZN(n1998) );
  aoi22d1 U2643 ( .A1(\RegFilePlugin_regFile[10][2] ), .A2(n1993), .B1(
        \RegFilePlugin_regFile[23][2] ), .B2(n1544), .ZN(n1997) );
  aoi22d1 U2644 ( .A1(\RegFilePlugin_regFile[25][2] ), .A2(n1607), .B1(
        \RegFilePlugin_regFile[18][2] ), .B2(n1952), .ZN(n1996) );
  aoi22d1 U2645 ( .A1(\RegFilePlugin_regFile[26][2] ), .A2(n1649), .B1(
        \RegFilePlugin_regFile[15][2] ), .B2(n1994), .ZN(n1995) );
  or04d0 U2646 ( .A1(n2002), .A2(n2001), .A3(n2000), .A4(n1999), .Z(N885) );
  aoi22d1 U2647 ( .A1(\RegFilePlugin_regFile[4][4] ), .A2(n2004), .B1(
        \RegFilePlugin_regFile[14][4] ), .B2(n2003), .ZN(n2010) );
  aoi22d1 U2648 ( .A1(\RegFilePlugin_regFile[17][4] ), .A2(n2005), .B1(
        \RegFilePlugin_regFile[29][4] ), .B2(n1501), .ZN(n2009) );
  aoi22d1 U2649 ( .A1(\RegFilePlugin_regFile[20][4] ), .A2(n2006), .B1(
        \RegFilePlugin_regFile[25][4] ), .B2(n1607), .ZN(n2008) );
  aoi22d1 U2650 ( .A1(\RegFilePlugin_regFile[30][4] ), .A2(n1837), .B1(
        \RegFilePlugin_regFile[6][4] ), .B2(n1522), .ZN(n2007) );
  aoi22d1 U2651 ( .A1(\RegFilePlugin_regFile[16][4] ), .A2(n1671), .B1(
        \RegFilePlugin_regFile[9][4] ), .B2(n2011), .ZN(n2019) );
  aoi22d1 U2652 ( .A1(\RegFilePlugin_regFile[1][4] ), .A2(n2012), .B1(
        \RegFilePlugin_regFile[28][4] ), .B2(n1903), .ZN(n2018) );
  aoi22d1 U2653 ( .A1(\RegFilePlugin_regFile[11][4] ), .A2(n2013), .B1(
        \RegFilePlugin_regFile[21][4] ), .B2(n1377), .ZN(n2017) );
  aoi22d1 U2654 ( .A1(\RegFilePlugin_regFile[26][4] ), .A2(n2015), .B1(
        \RegFilePlugin_regFile[22][4] ), .B2(n2014), .ZN(n2016) );
  aoi22d1 U2655 ( .A1(\RegFilePlugin_regFile[23][4] ), .A2(n2021), .B1(
        \RegFilePlugin_regFile[24][4] ), .B2(n2020), .ZN(n2029) );
  aoi22d1 U2656 ( .A1(\RegFilePlugin_regFile[5][4] ), .A2(n1606), .B1(
        \RegFilePlugin_regFile[3][4] ), .B2(n2022), .ZN(n2028) );
  aoi22d1 U2657 ( .A1(\RegFilePlugin_regFile[7][4] ), .A2(n1543), .B1(
        \RegFilePlugin_regFile[15][4] ), .B2(n2023), .ZN(n2027) );
  aoi22d1 U2658 ( .A1(\RegFilePlugin_regFile[13][4] ), .A2(n2025), .B1(
        \RegFilePlugin_regFile[19][4] ), .B2(n2024), .ZN(n2026) );
  aoi22d1 U2659 ( .A1(\RegFilePlugin_regFile[0][4] ), .A2(n2030), .B1(
        \RegFilePlugin_regFile[18][4] ), .B2(n1952), .ZN(n2037) );
  aoi22d1 U2660 ( .A1(\RegFilePlugin_regFile[10][4] ), .A2(n1416), .B1(
        \RegFilePlugin_regFile[8][4] ), .B2(n1670), .ZN(n2036) );
  aoi22d1 U2661 ( .A1(\RegFilePlugin_regFile[2][4] ), .A2(n2032), .B1(
        \RegFilePlugin_regFile[12][4] ), .B2(n2031), .ZN(n2035) );
  aoi22d1 U2662 ( .A1(\RegFilePlugin_regFile[27][4] ), .A2(n2033), .B1(
        \RegFilePlugin_regFile[31][4] ), .B2(n1417), .ZN(n2034) );
  or04d0 U2663 ( .A1(n2041), .A2(n2040), .A3(n2039), .A4(n2038), .Z(N883) );
  nr02d0 U2664 ( .A1(writeBack_MEMORY_ADDRESS_LOW[1]), .A2(
        writeBack_MEMORY_ADDRESS_LOW[0]), .ZN(n2462) );
  inv0d0 U2665 ( .I(writeBack_MEMORY_ADDRESS_LOW[1]), .ZN(n2042) );
  an02d0 U2666 ( .A1(n2042), .A2(writeBack_MEMORY_ADDRESS_LOW[0]), .Z(n2458)
         );
  aoi22d1 U2667 ( .A1(n2462), .A2(iBus_rsp_payload_data[1]), .B1(n2458), .B2(
        iBus_rsp_payload_data[9]), .ZN(n2045) );
  nd02d0 U2668 ( .A1(writeBack_MEMORY_ADDRESS_LOW[1]), .A2(
        writeBack_MEMORY_ADDRESS_LOW[0]), .ZN(n2460) );
  inv0d0 U2669 ( .I(n2460), .ZN(n2453) );
  nr02d1 U2670 ( .A1(writeBack_MEMORY_ADDRESS_LOW[0]), .A2(n2042), .ZN(n2483)
         );
  aoi22d1 U2671 ( .A1(n2453), .A2(iBus_rsp_payload_data[25]), .B1(n2483), .B2(
        iBus_rsp_payload_data[17]), .ZN(n2044) );
  an02d0 U2672 ( .A1(lastStageIsValid), .A2(writeBack_MEMORY_ENABLE), .Z(n2476) );
  nd02d0 U2673 ( .A1(n2526), .A2(writeBack_REGFILE_WRITE_DATA[1]), .ZN(n2043)
         );
  aon211d1 U2674 ( .C1(n2045), .C2(n2044), .B(n2526), .A(n2043), .ZN(n3285) );
  inv0d0 U2675 ( .I(n3285), .ZN(n3429) );
  inv0d2 U2676 ( .I(n2428), .ZN(n2530) );
  nd02d4 U2677 ( .A1(lastStageIsValid), .A2(n2530), .ZN(n2531) );
  nd02d1 U2678 ( .A1(n2530), .A2(n2046), .ZN(n2514) );
  inv0d0 U2679 ( .I(DebugPlugin_busReadDataReg[1]), .ZN(n2059) );
  oai22d1 U2680 ( .A1(n3429), .A2(n2531), .B1(n2514), .B2(n2059), .ZN(n6071)
         );
  aoi22d1 U2681 ( .A1(n2462), .A2(iBus_rsp_payload_data[0]), .B1(n2458), .B2(
        iBus_rsp_payload_data[8]), .ZN(n2049) );
  aoi22d1 U2682 ( .A1(n2453), .A2(iBus_rsp_payload_data[24]), .B1(n2483), .B2(
        iBus_rsp_payload_data[16]), .ZN(n2048) );
  nd02d0 U2683 ( .A1(n2526), .A2(writeBack_REGFILE_WRITE_DATA[0]), .ZN(n2047)
         );
  aon211d1 U2684 ( .C1(n2049), .C2(n2048), .B(n2526), .A(n2047), .ZN(n3251) );
  inv0d0 U2685 ( .I(n3251), .ZN(n3394) );
  inv0d0 U2686 ( .I(DebugPlugin_busReadDataReg[0]), .ZN(n2058) );
  oai22d1 U2687 ( .A1(n3394), .A2(n2531), .B1(n2514), .B2(n2058), .ZN(n6072)
         );
  inv0d0 U2688 ( .I(CsrPlugin_exceptionPortCtrl_exceptionContext_code[0]), 
        .ZN(n3670) );
  oai21d1 U2689 ( .B1(n2134), .B2(n3670), .A(n2193), .ZN(n6211) );
  inv0d0 U2690 ( .I(n3672), .ZN(n3677) );
  aor22d1 U2691 ( .A1(CsrPlugin_hadException), .A2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_code[2]), .B1(n3677), 
        .B2(CsrPlugin_mcause_exceptionCode[2]), .Z(n4075) );
  nd03d0 U2692 ( .A1(CsrPlugin_mstatus_MIE), .A2(CsrPlugin_mie_MSIE), .A3(
        CsrPlugin_mip_MSIP), .ZN(n3669) );
  nd03d0 U2693 ( .A1(CsrPlugin_mip_MEIP), .A2(CsrPlugin_mie_MEIE), .A3(
        CsrPlugin_mstatus_MIE), .ZN(n3668) );
  inv0d0 U2694 ( .I(n2534), .ZN(n3675) );
  aoi211d1 U2695 ( .C1(n3669), .C2(n3668), .A(n3675), .B(reset), .ZN(N1785) );
  oai21d1 U2696 ( .B1(CsrPlugin_exceptionPendings_1), .B2(n2051), .A(n2050), 
        .ZN(n2369) );
  nd02d0 U2697 ( .A1(n7121), .A2(n2589), .ZN(n2052) );
  oai22d1 U2698 ( .A1(n2362), .A2(n2240), .B1(n2369), .B2(n2052), .ZN(N1783)
         );
  inv0d2 U2699 ( .I(n2621), .ZN(n3558) );
  nd02d0 U2700 ( .A1(n3818), .A2(n2368), .ZN(n2055) );
  oan211d1 U2701 ( .C1(n3558), .C2(n2369), .B(n2055), .A(n2412), .ZN(N1782) );
  nr02d0 U2702 ( .A1(switch_Fetcher_l362[1]), .A2(switch_Fetcher_l362[0]), 
        .ZN(n2235) );
  nr04d0 U2703 ( .A1(debug_bus_cmd_payload_address[5]), .A2(
        debug_bus_cmd_payload_address[4]), .A3(
        debug_bus_cmd_payload_address[3]), .A4(
        debug_bus_cmd_payload_address[7]), .ZN(n2056) );
  nd03d0 U2704 ( .A1(n2056), .A2(debug_bus_cmd_payload_wr), .A3(
        debug_bus_cmd_valid), .ZN(n2057) );
  nr02d0 U2705 ( .A1(n2057), .A2(debug_bus_cmd_payload_address[6]), .ZN(n2415)
         );
  nd02d0 U2706 ( .A1(debug_bus_cmd_payload_address[2]), .A2(n2415), .ZN(n2228)
         );
  aor21d1 U2707 ( .B1(switch_Fetcher_l362[2]), .B2(n2235), .A(n2228), .Z(
        debug_bus_cmd_ready) );
  aoim22d1 U2708 ( .A1(_zz_when_DebugPlugin_l244), .A2(n2058), .B1(
        DebugPlugin_resetIt), .B2(_zz_when_DebugPlugin_l244), .Z(
        debug_bus_rsp_data[0]) );
  aoi22d1 U2709 ( .A1(_zz_when_DebugPlugin_l244), .A2(n2059), .B1(n2435), .B2(
        n7264), .ZN(debug_bus_rsp_data[1]) );
  inv0d0 U2710 ( .I(DebugPlugin_busReadDataReg[2]), .ZN(n2440) );
  aoim22d1 U2711 ( .A1(_zz_when_DebugPlugin_l244), .A2(n2440), .B1(
        DebugPlugin_isPipBusy), .B2(_zz_when_DebugPlugin_l244), .Z(
        debug_bus_rsp_data[2]) );
  inv0d0 U2712 ( .I(DebugPlugin_busReadDataReg[3]), .ZN(n2444) );
  inv0d0 U2713 ( .I(DebugPlugin_haltedByBreak), .ZN(n2418) );
  aoi22d1 U2714 ( .A1(_zz_when_DebugPlugin_l244), .A2(n2444), .B1(n2418), .B2(
        n7264), .ZN(debug_bus_rsp_data[3]) );
  inv0d0 U2715 ( .I(DebugPlugin_busReadDataReg[4]), .ZN(n2448) );
  aoi22d1 U2716 ( .A1(_zz_when_DebugPlugin_l244), .A2(n2448), .B1(n2422), .B2(
        n7264), .ZN(debug_bus_rsp_data[4]) );
  inv0d0 U2717 ( .I(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[0] ), 
        .ZN(n3097) );
  nd03d0 U2718 ( .A1(iBus_rsp_valid), .A2(\iBusWishbone_ADR[3]_BAR ), .A3(
        n3097), .ZN(n3158) );
  nr03d0 U2719 ( .A1(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[1] ), 
        .A2(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[2] ), 
        .A3(n3158), .ZN(n3191) );
  buffd1 U2720 ( .I(n3191), .Z(n3197) );
  buffd1 U2721 ( .I(n3191), .Z(n3207) );
  aoim22d1 U2722 ( .A1(n3197), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[0][31] ), .B2(n3207), .Z(n6246) );
  inv0d0 U2723 ( .I(\IBusCachedPlugin_cache/n23 ), .ZN(n5321) );
  nr02d1 U2724 ( .A1(n3052), .A2(n2374), .ZN(n2356) );
  inv0d0 U2725 ( .I(n6936), .ZN(n7007) );
  nr03d0 U2726 ( .A1(switch_Fetcher_l362[2]), .A2(switch_Fetcher_l362[1]), 
        .A3(switch_Fetcher_l362[0]), .ZN(n2079) );
  buffd1 U2727 ( .I(n2079), .Z(n2086) );
  nd02d1 U2728 ( .A1(n7007), .A2(n2086), .ZN(n2097) );
  buffd1 U2729 ( .I(n2097), .Z(n2092) );
  aoi22d1 U2730 ( .A1(n2095), .A2(_zz_decode_LEGAL_INSTRUCTION_1[0]), .B1(
        debug_bus_cmd_payload_data[0]), .B2(n2094), .ZN(n2060) );
  oai21d1 U2731 ( .B1(n5321), .B2(n2092), .A(n2060), .ZN(n6245) );
  inv0d0 U2732 ( .I(\IBusCachedPlugin_cache/n22 ), .ZN(n7111) );
  aoi22d1 U2733 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[1]), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[1]), .B2(n2094), .ZN(n2061) );
  oai21d1 U2734 ( .B1(n7111), .B2(n2092), .A(n2061), .ZN(n6244) );
  inv0d0 U2735 ( .I(\IBusCachedPlugin_cache/n21 ), .ZN(n6255) );
  aoi22d1 U2736 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[2]), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[2]), .B2(n2094), .ZN(n2062) );
  oai21d1 U2737 ( .B1(n6255), .B2(n2092), .A(n2062), .ZN(n6243) );
  inv0d0 U2738 ( .I(\IBusCachedPlugin_cache/n20 ), .ZN(n6433) );
  aoi22d1 U2739 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[3]), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[3]), .B2(n2094), .ZN(n2063) );
  oai21d1 U2740 ( .B1(n6433), .B2(n2092), .A(n2063), .ZN(n6242) );
  inv0d0 U2741 ( .I(\IBusCachedPlugin_cache/n19 ), .ZN(n6799) );
  inv0d0 U2742 ( .I(debug_bus_cmd_payload_data[4]), .ZN(n2424) );
  inv0d1 U2743 ( .I(n2095), .ZN(n2088) );
  oai222d1 U2744 ( .A1(n2097), .A2(n6799), .B1(n2424), .B2(n2079), .C1(n2553), 
        .C2(n2088), .ZN(n6241) );
  inv0d0 U2745 ( .I(\IBusCachedPlugin_cache/n18 ), .ZN(n6780) );
  aoi22d1 U2746 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[5]), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[5]), .B2(n2094), .ZN(n2064) );
  oai21d1 U2747 ( .B1(n6780), .B2(n2092), .A(n2064), .ZN(n6240) );
  inv0d0 U2748 ( .I(\IBusCachedPlugin_cache/n17 ), .ZN(n6766) );
  aoi22d1 U2749 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[6]), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[6]), .B2(n2094), .ZN(n2065) );
  oai21d1 U2750 ( .B1(n6766), .B2(n2092), .A(n2065), .ZN(n6239) );
  inv0d0 U2751 ( .I(\IBusCachedPlugin_cache/n16 ), .ZN(n6752) );
  aoi22d1 U2752 ( .A1(decode_INSTRUCTION_7), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[7]), .B2(n2094), .ZN(n2066) );
  oai21d1 U2753 ( .B1(n6752), .B2(n2097), .A(n2066), .ZN(n6238) );
  inv0d0 U2754 ( .I(\IBusCachedPlugin_cache/n15 ), .ZN(n6737) );
  aoi22d1 U2755 ( .A1(decode_INSTRUCTION_8), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[8]), .B2(n2094), .ZN(n2067) );
  oai21d1 U2756 ( .B1(n6737), .B2(n2097), .A(n2067), .ZN(n6237) );
  inv0d0 U2757 ( .I(\IBusCachedPlugin_cache/n14 ), .ZN(n6721) );
  aoi22d1 U2758 ( .A1(decode_INSTRUCTION_9), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[9]), .B2(n2094), .ZN(n2068) );
  oai21d1 U2759 ( .B1(n6721), .B2(n2092), .A(n2068), .ZN(n6236) );
  inv0d0 U2760 ( .I(\IBusCachedPlugin_cache/n13 ), .ZN(n6708) );
  aoi22d1 U2761 ( .A1(decode_INSTRUCTION_10), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[10]), .B2(n2094), .ZN(n2069) );
  oai21d1 U2762 ( .B1(n6708), .B2(n2097), .A(n2069), .ZN(n6235) );
  inv0d0 U2763 ( .I(\IBusCachedPlugin_cache/n12 ), .ZN(n6693) );
  aoi22d1 U2764 ( .A1(decode_INSTRUCTION_11), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[11]), .B2(n2094), .ZN(n2070) );
  oai21d1 U2765 ( .B1(n6693), .B2(n2097), .A(n2070), .ZN(n6234) );
  inv0d0 U2766 ( .I(\IBusCachedPlugin_cache/n11 ), .ZN(n6680) );
  inv0d0 U2767 ( .I(debug_bus_cmd_payload_data[12]), .ZN(n2071) );
  oai222d1 U2768 ( .A1(n2092), .A2(n6680), .B1(n2071), .B2(n2079), .C1(n2554), 
        .C2(n2088), .ZN(n6233) );
  inv0d0 U2769 ( .I(\IBusCachedPlugin_cache/n10 ), .ZN(n6664) );
  inv0d0 U2770 ( .I(debug_bus_cmd_payload_data[13]), .ZN(n2073) );
  oai222d1 U2771 ( .A1(n2097), .A2(n6664), .B1(n2073), .B2(n2079), .C1(n2072), 
        .C2(n2088), .ZN(n6232) );
  inv0d0 U2772 ( .I(\IBusCachedPlugin_cache/n9 ), .ZN(n6649) );
  aoi22d1 U2773 ( .A1(\_zz_decode_LEGAL_INSTRUCTION_7[14] ), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[14]), .B2(n2094), .ZN(n2074) );
  oai21d1 U2774 ( .B1(n6649), .B2(n2097), .A(n2074), .ZN(n6231) );
  inv0d0 U2775 ( .I(debug_bus_cmd_payload_data[15]), .ZN(n2075) );
  oai222d1 U2776 ( .A1(n2092), .A2(n6636), .B1(n2075), .B2(n2079), .C1(n174), 
        .C2(n2088), .ZN(n6230) );
  inv0d0 U2777 ( .I(IBusCachedPlugin_cache_io_cpu_fetch_data[16]), .ZN(n6623)
         );
  inv0d0 U2778 ( .I(debug_bus_cmd_payload_data[16]), .ZN(n2076) );
  oai222d1 U2779 ( .A1(n2097), .A2(n6623), .B1(n2076), .B2(n2079), .C1(n2623), 
        .C2(n2088), .ZN(n6229) );
  inv0d0 U2780 ( .I(debug_bus_cmd_payload_data[17]), .ZN(n2077) );
  oai222d1 U2781 ( .A1(n2092), .A2(n6611), .B1(n2077), .B2(n2079), .C1(n2622), 
        .C2(n2088), .ZN(n6228) );
  inv0d0 U2782 ( .I(debug_bus_cmd_payload_data[18]), .ZN(n2078) );
  oai222d1 U2783 ( .A1(n2092), .A2(n6598), .B1(n2078), .B2(n2079), .C1(n173), 
        .C2(n2088), .ZN(n6227) );
  inv0d0 U2784 ( .I(debug_bus_cmd_payload_data[19]), .ZN(n2080) );
  oai222d1 U2785 ( .A1(n2097), .A2(n6586), .B1(n2080), .B2(n2079), .C1(n2618), 
        .C2(n2088), .ZN(n6226) );
  inv0d0 U2786 ( .I(IBusCachedPlugin_cache_io_cpu_fetch_data[20]), .ZN(n6574)
         );
  inv0d0 U2787 ( .I(debug_bus_cmd_payload_data[20]), .ZN(n2081) );
  oai222d1 U2788 ( .A1(n2092), .A2(n6574), .B1(n2081), .B2(n2086), .C1(n2617), 
        .C2(n2088), .ZN(n6225) );
  inv0d0 U2789 ( .I(debug_bus_cmd_payload_data[21]), .ZN(n2082) );
  oai222d1 U2790 ( .A1(n2097), .A2(n6562), .B1(n2082), .B2(n2086), .C1(n2616), 
        .C2(n2088), .ZN(n6224) );
  inv0d0 U2791 ( .I(IBusCachedPlugin_cache_io_cpu_fetch_data[22]), .ZN(n6549)
         );
  inv0d0 U2792 ( .I(debug_bus_cmd_payload_data[22]), .ZN(n2083) );
  oai222d1 U2793 ( .A1(n2097), .A2(n6549), .B1(n2083), .B2(n2086), .C1(n2615), 
        .C2(n2088), .ZN(n6223) );
  inv0d0 U2794 ( .I(IBusCachedPlugin_cache_io_cpu_fetch_data[23]), .ZN(n6536)
         );
  inv0d0 U2795 ( .I(debug_bus_cmd_payload_data[23]), .ZN(n2084) );
  oai222d1 U2796 ( .A1(n2097), .A2(n6536), .B1(n2084), .B2(n2086), .C1(n2614), 
        .C2(n2088), .ZN(n6222) );
  inv0d0 U2797 ( .I(debug_bus_cmd_payload_data[24]), .ZN(n2085) );
  oai222d1 U2798 ( .A1(n2097), .A2(n6523), .B1(n2085), .B2(n2086), .C1(n2613), 
        .C2(n2088), .ZN(n6221) );
  inv0d0 U2799 ( .I(debug_bus_cmd_payload_data[25]), .ZN(n2420) );
  inv0d0 U2800 ( .I(\IBusCachedPlugin_cache/n8 ), .ZN(n6511) );
  oai222d1 U2801 ( .A1(n2612), .A2(n2088), .B1(n2420), .B2(n2086), .C1(n6511), 
        .C2(n2092), .ZN(n6220) );
  inv0d0 U2802 ( .I(debug_bus_cmd_payload_data[26]), .ZN(n2087) );
  inv0d0 U2803 ( .I(\IBusCachedPlugin_cache/n7 ), .ZN(n6499) );
  oai222d1 U2804 ( .A1(n2610), .A2(n2088), .B1(n2087), .B2(n2086), .C1(n6499), 
        .C2(n2092), .ZN(n6219) );
  inv0d0 U2805 ( .I(\IBusCachedPlugin_cache/n6 ), .ZN(n6487) );
  aoi22d1 U2806 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13[27]), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[27]), .B2(n2094), .ZN(n2089) );
  oai21d1 U2807 ( .B1(n6487), .B2(n2092), .A(n2089), .ZN(n6218) );
  inv0d0 U2808 ( .I(\IBusCachedPlugin_cache/n5 ), .ZN(n6473) );
  aoi22d1 U2809 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13[28]), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[28]), .B2(n2094), .ZN(n2090) );
  oai21d1 U2810 ( .B1(n6473), .B2(n2092), .A(n2090), .ZN(n6217) );
  inv0d0 U2811 ( .I(\IBusCachedPlugin_cache/n4 ), .ZN(n6458) );
  aoi22d1 U2812 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13[29]), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[29]), .B2(n2094), .ZN(n2091) );
  oai21d1 U2813 ( .B1(n6458), .B2(n2092), .A(n2091), .ZN(n6216) );
  inv0d0 U2814 ( .I(\IBusCachedPlugin_cache/n3 ), .ZN(n6446) );
  aoi22d1 U2815 ( .A1(decode_INSTRUCTION_30), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[30]), .B2(n2094), .ZN(n2093) );
  oai21d1 U2816 ( .B1(n6446), .B2(n2097), .A(n2093), .ZN(n6215) );
  inv0d0 U2817 ( .I(\IBusCachedPlugin_cache/n2 ), .ZN(n3733) );
  aoi22d1 U2818 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13_31), .A2(n2095), .B1(
        debug_bus_cmd_payload_data[31]), .B2(n2094), .ZN(n2096) );
  oai21d1 U2819 ( .B1(n3733), .B2(n2097), .A(n2096), .ZN(n6214) );
  nr03d0 U2820 ( .A1(\_zz__zz_decode_ENV_CTRL_2_1[20] ), .A2(
        decode_INSTRUCTION_21), .A3(n2610), .ZN(n2548) );
  inv0d0 U2821 ( .I(_zz_decode_LEGAL_INSTRUCTION_13[27]), .ZN(n2608) );
  inv0d0 U2822 ( .I(_zz_decode_LEGAL_INSTRUCTION_13_31), .ZN(n2603) );
  nr04d0 U2823 ( .A1(n3238), .A2(n2608), .A3(n2603), .A4(n2098), .ZN(n2099) );
  nd04d0 U2824 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13[29]), .A2(n2559), .A3(
        n2548), .A4(n2099), .ZN(n2536) );
  oai22d1 U2825 ( .A1(decode_INSTRUCTION_30), .A2(n2536), .B1(n3558), .B2(
        n2244), .ZN(n6213) );
  aoi22d1 U2826 ( .A1(n2109), .A2(execute_RS2[31]), .B1(n2105), .B2(
        execute_PC[31]), .ZN(n2100) );
  nd02d0 U2827 ( .A1(n2100), .A2(n305), .ZN(n2637) );
  inv0d0 U2828 ( .I(execute_RS1[30]), .ZN(n6257) );
  inv0d0 U2829 ( .I(_zz__zz_execute_SRC2_3[10]), .ZN(n2604) );
  oai22d1 U2830 ( .A1(n2111), .A2(n6257), .B1(n302), .B2(n2604), .ZN(n2659) );
  aoi22d1 U2831 ( .A1(n3026), .A2(n2637), .B1(n2969), .B2(n2659), .ZN(n2132)
         );
  inv0d0 U2832 ( .I(n2637), .ZN(n2123) );
  oai22d1 U2833 ( .A1(n2123), .A2(n2961), .B1(n2570), .B2(n314), .ZN(n2127) );
  inv0d0 U2834 ( .I(execute_RS1[31]), .ZN(n6256) );
  inv0d0 U2835 ( .I(n6343), .ZN(n6284) );
  oai22d1 U2836 ( .A1(n2111), .A2(n6256), .B1(n302), .B2(n6284), .ZN(n2649) );
  aoi22d1 U2837 ( .A1(n2123), .A2(n2110), .B1(n2117), .B2(n2637), .ZN(n2121)
         );
  aoi22d1 U2838 ( .A1(n2114), .A2(execute_RS2[30]), .B1(n2105), .B2(
        execute_PC[30]), .ZN(n2101) );
  nd02d0 U2839 ( .A1(n2101), .A2(n305), .ZN(n2658) );
  inv0d0 U2840 ( .I(n2658), .ZN(n2653) );
  aoi22d1 U2841 ( .A1(n2653), .A2(n2594), .B1(n2117), .B2(n2658), .ZN(n2651)
         );
  inv0d0 U2842 ( .I(execute_RS1[29]), .ZN(n6258) );
  inv0d0 U2843 ( .I(_zz__zz_execute_SRC2_3[9]), .ZN(n6459) );
  oai22d1 U2844 ( .A1(n2111), .A2(n6258), .B1(n302), .B2(n6459), .ZN(n2670) );
  aoi22d1 U2845 ( .A1(n2114), .A2(execute_RS2[29]), .B1(n2105), .B2(
        execute_PC[29]), .ZN(n2102) );
  nd02d0 U2846 ( .A1(n2102), .A2(n305), .ZN(n2665) );
  inv0d0 U2847 ( .I(n2665), .ZN(n2666) );
  aoi22d1 U2848 ( .A1(n2666), .A2(n2594), .B1(n2117), .B2(n2665), .ZN(n2668)
         );
  inv0d0 U2849 ( .I(execute_RS1[28]), .ZN(n6259) );
  inv0d0 U2850 ( .I(_zz__zz_execute_SRC2_3[8]), .ZN(n6474) );
  oai22d1 U2851 ( .A1(n2111), .A2(n6259), .B1(n302), .B2(n6474), .ZN(n2694) );
  aoi22d1 U2852 ( .A1(n2103), .A2(execute_RS2[28]), .B1(n2105), .B2(
        execute_PC[28]), .ZN(n2104) );
  nd02d0 U2853 ( .A1(n2104), .A2(n305), .ZN(n2689) );
  aoim22d1 U2854 ( .A1(n2117), .A2(n2689), .B1(n2689), .B2(n2117), .Z(n2680)
         );
  inv0d0 U2855 ( .I(execute_RS1[27]), .ZN(n6260) );
  inv0d0 U2856 ( .I(_zz__zz_execute_SRC2_3[7]), .ZN(n2607) );
  oai22d1 U2857 ( .A1(n2111), .A2(n6260), .B1(n302), .B2(n2607), .ZN(n2711) );
  aoi22d1 U2858 ( .A1(n2114), .A2(execute_RS2[27]), .B1(n2105), .B2(
        execute_PC[27]), .ZN(n2106) );
  nd02d0 U2859 ( .A1(n2106), .A2(n305), .ZN(n2695) );
  inv0d0 U2860 ( .I(n2695), .ZN(n2696) );
  aoi22d1 U2861 ( .A1(n2696), .A2(n2110), .B1(n2117), .B2(n2695), .ZN(n2699)
         );
  inv0d0 U2862 ( .I(execute_RS1[26]), .ZN(n6261) );
  inv0d0 U2863 ( .I(_zz__zz_execute_SRC2_3[6]), .ZN(n2609) );
  oai22d1 U2864 ( .A1(n2111), .A2(n6261), .B1(n302), .B2(n2609), .ZN(n2713) );
  aoi22d1 U2865 ( .A1(n2109), .A2(execute_RS2[26]), .B1(n2113), .B2(
        execute_PC[26]), .ZN(n2107) );
  nd02d0 U2866 ( .A1(n2107), .A2(n305), .ZN(n2712) );
  aoim22d1 U2867 ( .A1(n2117), .A2(n2712), .B1(n2712), .B2(n2117), .Z(n2709)
         );
  inv0d0 U2868 ( .I(execute_RS1[25]), .ZN(n6262) );
  inv0d0 U2869 ( .I(_zz__zz_execute_SRC2_3[5]), .ZN(n2611) );
  oai22d1 U2870 ( .A1(n2111), .A2(n6262), .B1(n302), .B2(n2611), .ZN(n2728) );
  oaim21d1 U2871 ( .B1(n2113), .B2(execute_PC[25]), .A(n305), .ZN(n2108) );
  aoi21d1 U2872 ( .B1(n2109), .B2(execute_RS2[25]), .A(n2108), .ZN(n2721) );
  inv0d0 U2873 ( .I(n2721), .ZN(n2722) );
  aoi22d1 U2874 ( .A1(n2721), .A2(n2110), .B1(n2117), .B2(n2722), .ZN(n2726)
         );
  inv0d0 U2875 ( .I(execute_RS1[24]), .ZN(n6263) );
  inv0d0 U2876 ( .I(_zz__zz_execute_BranchPlugin_branch_src2_3), .ZN(n6293) );
  oai22d1 U2877 ( .A1(n2111), .A2(n6263), .B1(n6293), .B2(n302), .ZN(n2740) );
  aoi22d1 U2878 ( .A1(n2114), .A2(execute_RS2[24]), .B1(n2113), .B2(
        execute_PC[24]), .ZN(n2112) );
  nd02d0 U2879 ( .A1(n2112), .A2(n305), .ZN(n2741) );
  aoim22d1 U2880 ( .A1(n2117), .A2(n2741), .B1(n2741), .B2(n2117), .Z(n2737)
         );
  aoi22d1 U2881 ( .A1(n2114), .A2(execute_RS2[23]), .B1(n2113), .B2(
        execute_PC[23]), .ZN(n2116) );
  nd02d0 U2882 ( .A1(n2116), .A2(n305), .ZN(n2759) );
  aoim22d1 U2883 ( .A1(n2117), .A2(n2759), .B1(n2759), .B2(n2117), .Z(n2757)
         );
  xr03d1 U2884 ( .A1(n2121), .A2(n2120), .A3(n2649), .Z(n2122) );
  aoi22d1 U2885 ( .A1(execute_SRC2_FORCE_ZERO), .A2(n2649), .B1(n2122), .B2(
        n2897), .ZN(n6805) );
  nd02d0 U2886 ( .A1(n2123), .A2(n2649), .ZN(n2633) );
  oai21d1 U2887 ( .B1(n2123), .B2(n2649), .A(n2633), .ZN(n3754) );
  aoi22d1 U2888 ( .A1(n3029), .A2(memory_REGFILE_WRITE_DATA[30]), .B1(n2960), 
        .B2(n3754), .ZN(n2125) );
  nd03d0 U2889 ( .A1(execute_SHIFT_CTRL[0]), .A2(n2818), .A3(
        memory_REGFILE_WRITE_DATA[31]), .ZN(n2124) );
  oai211d1 U2890 ( .C1(n6805), .C2(n3005), .A(n2125), .B(n2124), .ZN(n2126) );
  oan211d1 U2891 ( .C1(n3026), .C2(n2127), .B(n2649), .A(n2126), .ZN(n2131) );
  aoi22d1 U2892 ( .A1(CsrPlugin_mepc[31]), .A2(execute_CsrPlugin_csr_833), 
        .B1(CsrPlugin_mtval[31]), .B2(n2327), .ZN(n2129) );
  aoi22d1 U2893 ( .A1(CsrPlugin_mcause_interrupt), .A2(
        execute_CsrPlugin_csr_834), .B1(
        _zz_CsrPlugin_csrMapping_readDataInit[31]), .B2(n2328), .ZN(n2128) );
  nd02d0 U2894 ( .A1(n2129), .A2(n2128), .ZN(n2249) );
  aoi22d1 U2895 ( .A1(n2999), .A2(n2249), .B1(memory_REGFILE_WRITE_DATA[31]), 
        .B2(n299), .ZN(n2130) );
  aon211d1 U2896 ( .C1(n2132), .C2(n2131), .B(n2996), .A(n2130), .ZN(n6212) );
  inv0d0 U2897 ( .I(CsrPlugin_exceptionPortCtrl_exceptionContext_code[3]), 
        .ZN(n2133) );
  oai21d1 U2898 ( .B1(n2134), .B2(n2133), .A(n2189), .ZN(n6210) );
  oaim21d1 U2899 ( .B1(n2204), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_code[2]), .A(n2135), .ZN(
        n6209) );
  aoi22d1 U2900 ( .A1(memory_BRANCH_CALC[31]), .A2(n2150), .B1(
        memory_REGFILE_WRITE_DATA[31]), .B2(n2198), .ZN(n2139) );
  aoi22d1 U2901 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13_31), .A2(n2186), .B1(
        n2204), .B2(CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[31]), 
        .ZN(n2138) );
  oai211d1 U2902 ( .C1(n6284), .C2(n2193), .A(n2139), .B(n2138), .ZN(n6206) );
  buffd1 U2903 ( .I(n2150), .Z(n2203) );
  aoi22d1 U2904 ( .A1(memory_BRANCH_CALC[30]), .A2(n2203), .B1(
        memory_REGFILE_WRITE_DATA[30]), .B2(n2198), .ZN(n2141) );
  aoi22d1 U2905 ( .A1(decode_INSTRUCTION_30), .A2(n2186), .B1(n2204), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[30]), .ZN(n2140)
         );
  oai211d1 U2906 ( .C1(n2604), .C2(n2193), .A(n2141), .B(n2140), .ZN(n6205) );
  aoi22d1 U2907 ( .A1(memory_BRANCH_CALC[29]), .A2(n2150), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[29]), .ZN(n2143) );
  aoi22d1 U2908 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13[29]), .A2(n2186), .B1(
        n2204), .B2(CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[29]), 
        .ZN(n2142) );
  oai211d1 U2909 ( .C1(n6459), .C2(n2193), .A(n2143), .B(n2142), .ZN(n6204) );
  aoi22d1 U2910 ( .A1(memory_BRANCH_CALC[28]), .A2(n2203), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[28]), .ZN(n2145) );
  aoi22d1 U2911 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13[28]), .A2(n2186), .B1(
        n2204), .B2(CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[28]), 
        .ZN(n2144) );
  oai211d1 U2912 ( .C1(n6474), .C2(n2193), .A(n2145), .B(n2144), .ZN(n6203) );
  buffd1 U2913 ( .I(n2150), .Z(n2207) );
  aoi22d1 U2914 ( .A1(memory_BRANCH_CALC[27]), .A2(n2207), .B1(
        memory_REGFILE_WRITE_DATA[27]), .B2(n2198), .ZN(n2147) );
  aoi22d1 U2915 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13[27]), .A2(n2186), .B1(
        n2204), .B2(CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[27]), 
        .ZN(n2146) );
  oai211d1 U2916 ( .C1(n2607), .C2(n2193), .A(n2147), .B(n2146), .ZN(n6202) );
  aoi22d1 U2917 ( .A1(memory_BRANCH_CALC[26]), .A2(n2150), .B1(
        memory_REGFILE_WRITE_DATA[26]), .B2(n2198), .ZN(n2149) );
  buffd1 U2918 ( .I(n2181), .Z(n2208) );
  aoi22d1 U2919 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13[26]), .A2(n2186), .B1(
        n2208), .B2(CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[26]), 
        .ZN(n2148) );
  oai211d1 U2920 ( .C1(n2609), .C2(n2193), .A(n2149), .B(n2148), .ZN(n6201) );
  aoi22d1 U2921 ( .A1(memory_BRANCH_CALC[25]), .A2(n2150), .B1(
        memory_REGFILE_WRITE_DATA[25]), .B2(n2198), .ZN(n2152) );
  aoi22d1 U2922 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13[25]), .A2(n2190), .B1(
        n2208), .B2(CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[25]), 
        .ZN(n2151) );
  oai211d1 U2923 ( .C1(n2611), .C2(n2189), .A(n2152), .B(n2151), .ZN(n6200) );
  aoi22d1 U2924 ( .A1(memory_BRANCH_CALC[24]), .A2(n2207), .B1(
        memory_REGFILE_WRITE_DATA[24]), .B2(n2198), .ZN(n2154) );
  aoi22d1 U2925 ( .A1(decode_INSTRUCTION_24), .A2(n2186), .B1(n2208), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[24]), .ZN(n2153)
         );
  oai211d1 U2926 ( .C1(n6293), .C2(n2193), .A(n2154), .B(n2153), .ZN(n6199) );
  aoi22d1 U2927 ( .A1(memory_BRANCH_CALC[23]), .A2(n2207), .B1(
        memory_REGFILE_WRITE_DATA[23]), .B2(n2198), .ZN(n2156) );
  aoi22d1 U2928 ( .A1(decode_INSTRUCTION_23), .A2(n2190), .B1(n2208), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[23]), .ZN(n2155)
         );
  oai211d1 U2929 ( .C1(n6295), .C2(n2189), .A(n2156), .B(n2155), .ZN(n6198) );
  aoi22d1 U2930 ( .A1(memory_BRANCH_CALC[22]), .A2(n2207), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[22]), .ZN(n2158) );
  aoi22d1 U2931 ( .A1(decode_INSTRUCTION_22), .A2(n2186), .B1(n2208), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[22]), .ZN(n2157)
         );
  oai211d1 U2932 ( .C1(n6298), .C2(n2193), .A(n2158), .B(n2157), .ZN(n6197) );
  aoi22d1 U2933 ( .A1(memory_BRANCH_CALC[21]), .A2(n2207), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[21]), .ZN(n2160) );
  aoi22d1 U2934 ( .A1(decode_INSTRUCTION_21), .A2(n2190), .B1(n2208), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[21]), .ZN(n2159)
         );
  oai211d1 U2935 ( .C1(n6303), .C2(n2189), .A(n2160), .B(n2159), .ZN(n6196) );
  aoi22d1 U2936 ( .A1(memory_BRANCH_CALC[20]), .A2(n2207), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[20]), .ZN(n2162) );
  aoi22d1 U2937 ( .A1(\_zz__zz_decode_ENV_CTRL_2_1[20] ), .A2(n2186), .B1(
        n2208), .B2(CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[20]), 
        .ZN(n2161) );
  oai211d1 U2938 ( .C1(n6307), .C2(n2193), .A(n2162), .B(n2161), .ZN(n6195) );
  aoi22d1 U2939 ( .A1(memory_BRANCH_CALC[19]), .A2(n2207), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[19]), .ZN(n2164) );
  aoi22d1 U2940 ( .A1(decode_INSTRUCTION[19]), .A2(n2190), .B1(n2208), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[19]), .ZN(n2163)
         );
  oai211d1 U2941 ( .C1(n6269), .C2(n2189), .A(n2164), .B(n2163), .ZN(n6194) );
  aoi22d1 U2942 ( .A1(memory_BRANCH_CALC[18]), .A2(n2207), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[18]), .ZN(n2166) );
  aoi22d1 U2943 ( .A1(decode_INSTRUCTION[18]), .A2(n2186), .B1(n2208), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[18]), .ZN(n2165)
         );
  oai211d1 U2944 ( .C1(n6271), .C2(n2189), .A(n2166), .B(n2165), .ZN(n6193) );
  inv0d1 U2945 ( .I(n2186), .ZN(n2212) );
  aoi22d1 U2946 ( .A1(memory_BRANCH_CALC[17]), .A2(n2207), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[17]), .ZN(n2168) );
  aoi22d1 U2947 ( .A1(_zz__zz_execute_SRC1_1[2]), .A2(n2209), .B1(n2204), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[17]), .ZN(n2167)
         );
  oai211d1 U2948 ( .C1(n2622), .C2(n2212), .A(n2168), .B(n2167), .ZN(n6192) );
  aoi22d1 U2949 ( .A1(memory_BRANCH_CALC[16]), .A2(n2207), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[16]), .ZN(n2170) );
  aoi22d1 U2950 ( .A1(_zz__zz_execute_SRC1_1[1]), .A2(n2209), .B1(n2208), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[16]), .ZN(n2169)
         );
  oai211d1 U2951 ( .C1(n2623), .C2(n2212), .A(n2170), .B(n2169), .ZN(n6191) );
  aoi22d1 U2952 ( .A1(memory_BRANCH_CALC[15]), .A2(n2207), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[15]), .ZN(n2172) );
  aoi22d1 U2953 ( .A1(_zz__zz_execute_SRC1_1[0]), .A2(n2209), .B1(n2208), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[15]), .ZN(n2171)
         );
  oai211d1 U2954 ( .C1(n174), .C2(n2212), .A(n2172), .B(n2171), .ZN(n6190) );
  aoi22d1 U2955 ( .A1(memory_BRANCH_CALC[14]), .A2(n2207), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[14]), .ZN(n2174) );
  aoi22d1 U2956 ( .A1(_zz__zz_execute_BranchPlugin_branch_src2[13]), .A2(n2209), .B1(n2204), .B2(CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[14]), 
        .ZN(n2173) );
  oai211d1 U2957 ( .C1(n2625), .C2(n2212), .A(n2174), .B(n2173), .ZN(n6189) );
  aoi22d1 U2958 ( .A1(memory_BRANCH_CALC[13]), .A2(n2203), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[13]), .ZN(n2176) );
  aoi22d1 U2959 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1_13), .A2(n2190), .B1(
        n2204), .B2(CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[13]), 
        .ZN(n2175) );
  oai211d1 U2960 ( .C1(n6666), .C2(n2189), .A(n2176), .B(n2175), .ZN(n6188) );
  aoi22d1 U2961 ( .A1(memory_BRANCH_CALC[12]), .A2(n2203), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[12]), .ZN(n2178) );
  aoi22d1 U2962 ( .A1(_zz_decode_LEGAL_INSTRUCTION_7_12), .A2(n2186), .B1(
        n2208), .B2(CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[12]), 
        .ZN(n2177) );
  oai211d1 U2963 ( .C1(n6681), .C2(n2193), .A(n2178), .B(n2177), .ZN(n6187) );
  aoi22d1 U2964 ( .A1(memory_BRANCH_CALC[11]), .A2(n2203), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[11]), .ZN(n2180) );
  aoi22d1 U2965 ( .A1(_zz__zz_execute_SRC2_3[4]), .A2(n2209), .B1(n2208), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[11]), .ZN(n2179)
         );
  oai211d1 U2966 ( .C1(n2627), .C2(n2212), .A(n2180), .B(n2179), .ZN(n6186) );
  aoi22d1 U2967 ( .A1(memory_BRANCH_CALC[10]), .A2(n2203), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[10]), .ZN(n2183) );
  aoi22d1 U2968 ( .A1(_zz__zz_execute_SRC2_3[3]), .A2(n2209), .B1(n2181), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[10]), .ZN(n2182)
         );
  oai211d1 U2969 ( .C1(n2628), .C2(n2212), .A(n2183), .B(n2182), .ZN(n6185) );
  aoi22d1 U2970 ( .A1(memory_BRANCH_CALC[9]), .A2(n2203), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[9]), .ZN(n2185) );
  aoi22d1 U2971 ( .A1(decode_INSTRUCTION_9), .A2(n2186), .B1(n2204), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[9]), .ZN(n2184)
         );
  oai211d1 U2972 ( .C1(n6722), .C2(n2193), .A(n2185), .B(n2184), .ZN(n6184) );
  aoi22d1 U2973 ( .A1(memory_BRANCH_CALC[8]), .A2(n2203), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[8]), .ZN(n2188) );
  aoi22d1 U2974 ( .A1(decode_INSTRUCTION_8), .A2(n2186), .B1(n2204), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[8]), .ZN(n2187)
         );
  oai211d1 U2975 ( .C1(n6738), .C2(n2189), .A(n2188), .B(n2187), .ZN(n6183) );
  aoi22d1 U2976 ( .A1(memory_BRANCH_CALC[7]), .A2(n2203), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[7]), .ZN(n2192) );
  aoi22d1 U2977 ( .A1(decode_INSTRUCTION_7), .A2(n2190), .B1(n2208), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[7]), .ZN(n2191)
         );
  oai211d1 U2978 ( .C1(n6753), .C2(n2193), .A(n2192), .B(n2191), .ZN(n6182) );
  aoi22d1 U2979 ( .A1(memory_BRANCH_CALC[6]), .A2(n2203), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[6]), .ZN(n2195) );
  aoi22d1 U2980 ( .A1(n2209), .A2(execute_INSTRUCTION[6]), .B1(n2204), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[6]), .ZN(n2194)
         );
  oai211d1 U2981 ( .C1(n2577), .C2(n2212), .A(n2195), .B(n2194), .ZN(n6181) );
  aoi22d1 U2982 ( .A1(memory_BRANCH_CALC[5]), .A2(n2203), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[5]), .ZN(n2197) );
  aoi22d1 U2983 ( .A1(n2209), .A2(execute_INSTRUCTION[5]), .B1(n2208), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[5]), .ZN(n2196)
         );
  oai211d1 U2984 ( .C1(n2630), .C2(n2212), .A(n2197), .B(n2196), .ZN(n6180) );
  aoi22d1 U2985 ( .A1(memory_BRANCH_CALC[4]), .A2(n2203), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[4]), .ZN(n2200) );
  aoi22d1 U2986 ( .A1(n2209), .A2(execute_INSTRUCTION[4]), .B1(n2204), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[4]), .ZN(n2199)
         );
  oai211d1 U2987 ( .C1(n2553), .C2(n2212), .A(n2200), .B(n2199), .ZN(n6179) );
  aoi22d1 U2988 ( .A1(memory_BRANCH_CALC[3]), .A2(n2207), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[3]), .ZN(n2202) );
  aoi22d1 U2989 ( .A1(n2209), .A2(execute_INSTRUCTION[3]), .B1(n2204), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[3]), .ZN(n2201)
         );
  oai211d1 U2990 ( .C1(n2575), .C2(n2212), .A(n2202), .B(n2201), .ZN(n6178) );
  aoi22d1 U2991 ( .A1(memory_BRANCH_CALC[2]), .A2(n2203), .B1(n2198), .B2(
        memory_REGFILE_WRITE_DATA[2]), .ZN(n2206) );
  aoi22d1 U2992 ( .A1(n2209), .A2(execute_INSTRUCTION[2]), .B1(n2204), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[2]), .ZN(n2205)
         );
  oai211d1 U2993 ( .C1(n3047), .C2(n2212), .A(n2206), .B(n2205), .ZN(n6177) );
  inv0d0 U2994 ( .I(_zz_decode_LEGAL_INSTRUCTION_1[1]), .ZN(n3048) );
  aoi21d1 U2995 ( .B1(n2198), .B2(memory_REGFILE_WRITE_DATA[1]), .A(n2207), 
        .ZN(n2211) );
  aoi22d1 U2996 ( .A1(n2209), .A2(execute_INSTRUCTION[1]), .B1(n2208), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[1]), .ZN(n2210)
         );
  oai211d1 U2997 ( .C1(n3048), .C2(n2212), .A(n2211), .B(n2210), .ZN(n6176) );
  inv0d0 U2998 ( .I(n2213), .ZN(n2217) );
  aoi31d1 U2999 ( .B1(n2749), .B2(n2217), .B3(n2216), .A(n6977), .ZN(n2218) );
  aoi211d1 U3000 ( .C1(dBusWishbone_ACK), .C2(n7265), .A(n2412), .B(n2218), 
        .ZN(n6175) );
  inv0d0 U3001 ( .I(iBusWishbone_ADR[0]), .ZN(n2220) );
  an02d0 U3002 ( .A1(iBusWishbone_ACK), .A2(iBusWishbone_ADR[0]), .Z(n2224) );
  aoi211d1 U3003 ( .C1(n2220), .C2(n2219), .A(n2412), .B(n2224), .ZN(n6174) );
  nd02d0 U3004 ( .A1(n2224), .A2(iBusWishbone_ADR[1]), .ZN(n2221) );
  inv0d0 U3005 ( .I(n2221), .ZN(n2223) );
  inv0d0 U3006 ( .I(iBusWishbone_ADR[2]), .ZN(n2222) );
  aoi221d1 U3007 ( .B1(iBusWishbone_ADR[2]), .B2(n2223), .C1(n2222), .C2(n2221), .A(reset), .ZN(n6173) );
  aoim211d1 U3008 ( .C1(n2224), .C2(iBusWishbone_ADR[1]), .A(reset), .B(n2223), 
        .ZN(n6172) );
  inv0d0 U3009 ( .I(switch_Fetcher_l362[1]), .ZN(n2237) );
  nd02d0 U3010 ( .A1(n2234), .A2(n2237), .ZN(n2229) );
  aoi31d1 U3011 ( .B1(switch_Fetcher_l362[0]), .B2(n2234), .B3(n2237), .A(
        n2225), .ZN(n2238) );
  oai211d1 U3012 ( .C1(n2374), .C2(n2226), .A(n7121), .B(n2238), .ZN(n2236) );
  inv0d0 U3013 ( .I(n2236), .ZN(n2227) );
  oai21d1 U3014 ( .B1(n2229), .B2(n2228), .A(n2227), .ZN(n2232) );
  inv0d0 U3015 ( .I(switch_Fetcher_l362[0]), .ZN(n2231) );
  oai21d1 U3016 ( .B1(n2232), .B2(n2231), .A(n2230), .ZN(n6171) );
  nd03d0 U3017 ( .A1(switch_Fetcher_l362[0]), .A2(switch_Fetcher_l362[1]), 
        .A3(n2236), .ZN(n2233) );
  oan211d1 U3018 ( .C1(n2235), .C2(n2234), .B(n2233), .A(n2412), .ZN(n6170) );
  oai22d1 U3019 ( .A1(reset), .A2(n2238), .B1(n2237), .B2(n2236), .ZN(n6169)
         );
  nr13d1 U3020 ( .A1(memory_arbitration_isValid), .A2(n2241), .A3(n2239), .ZN(
        n6168) );
  nd02d0 U3021 ( .A1(execute_arbitration_isValid), .A2(n2358), .ZN(n2243) );
  oai22d1 U3022 ( .A1(n3235), .A2(n2243), .B1(n2241), .B2(n2240), .ZN(n6167)
         );
  inv0d1 U3023 ( .I(n3232), .ZN(n2620) );
  oai22d1 U3024 ( .A1(n2620), .A2(n2243), .B1(n2242), .B2(n2374), .ZN(n6166)
         );
  inv0d0 U3025 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[0]), .ZN(n2248) );
  inv0d0 U3026 ( .I(n3566), .ZN(n3561) );
  oai21d1 U3027 ( .B1(n2244), .B2(n3561), .A(n7121), .ZN(n2334) );
  inv0d0 U3028 ( .I(execute_CsrPlugin_csr_4032), .ZN(n2537) );
  aoi22d1 U3029 ( .A1(n2328), .A2(_zz_CsrPlugin_csrMapping_readDataInit[0]), 
        .B1(execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[0]), .ZN(n2246) );
  aoi22d1 U3030 ( .A1(execute_CsrPlugin_csr_834), .A2(
        CsrPlugin_mcause_exceptionCode[0]), .B1(execute_CsrPlugin_csr_833), 
        .B2(CsrPlugin_mepc[0]), .ZN(n2245) );
  oai211d1 U3031 ( .C1(n2537), .C2(n2247), .A(n2246), .B(n2245), .ZN(n2645) );
  inv0d0 U3032 ( .I(n2644), .ZN(n3036) );
  oai222d1 U3033 ( .A1(n2644), .A2(
        _zz__zz_execute_BranchPlugin_branch_src2[12]), .B1(n2644), .B2(n2645), 
        .C1(n3036), .C2(n2289), .ZN(n3568) );
  nd03d1 U3034 ( .A1(n2328), .A2(n3566), .A3(n7121), .ZN(n2322) );
  buffd1 U3035 ( .I(n2322), .Z(n2332) );
  oai22d1 U3036 ( .A1(n2248), .A2(n2334), .B1(n3568), .B2(n2332), .ZN(n6165)
         );
  inv0d0 U3037 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[31]), .ZN(n2250) );
  buffd1 U3038 ( .I(n2334), .Z(n2303) );
  inv0d0 U3039 ( .I(n2649), .ZN(n2638) );
  oai222d1 U3040 ( .A1(n2649), .A2(n2266), .B1(n2649), .B2(n2249), .C1(n2638), 
        .C2(n2289), .ZN(n3667) );
  oai22d1 U3041 ( .A1(n2250), .A2(n2303), .B1(n3667), .B2(n2332), .ZN(n6164)
         );
  inv0d0 U3042 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[30]), .ZN(n2252) );
  inv0d0 U3043 ( .I(CsrPlugin_mepc[30]), .ZN(n3658) );
  aoi22d1 U3044 ( .A1(execute_CsrPlugin_csr_3008), .A2(
        _zz_CsrPlugin_csrMapping_readDataInit[30]), .B1(
        execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[30]), .ZN(n2251) );
  oai21d1 U3045 ( .B1(n3658), .B2(n2541), .A(n2251), .ZN(n2660) );
  inv0d0 U3046 ( .I(n2659), .ZN(n2671) );
  oai222d1 U3047 ( .A1(n2659), .A2(n2266), .B1(n2659), .B2(n2660), .C1(n2671), 
        .C2(n2289), .ZN(n3661) );
  oai22d1 U3048 ( .A1(n2252), .A2(n2303), .B1(n3661), .B2(n2332), .ZN(n6163)
         );
  inv0d0 U3049 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[29]), .ZN(n2254) );
  inv0d0 U3050 ( .I(CsrPlugin_mepc[29]), .ZN(n3654) );
  aoi22d1 U3051 ( .A1(execute_CsrPlugin_csr_3008), .A2(
        _zz_CsrPlugin_csrMapping_readDataInit[29]), .B1(n2327), .B2(
        CsrPlugin_mtval[29]), .ZN(n2253) );
  oai21d1 U3052 ( .B1(n3654), .B2(n2541), .A(n2253), .ZN(n2664) );
  inv0d0 U3053 ( .I(n2670), .ZN(n2682) );
  oai222d1 U3054 ( .A1(n2670), .A2(n2266), .B1(n2670), .B2(n2664), .C1(n2682), 
        .C2(n2289), .ZN(n3655) );
  oai22d1 U3055 ( .A1(n2254), .A2(n2303), .B1(n3655), .B2(n2332), .ZN(n6162)
         );
  inv0d0 U3056 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[28]), .ZN(n2256) );
  inv0d0 U3057 ( .I(CsrPlugin_mepc[28]), .ZN(n3651) );
  aoi22d1 U3058 ( .A1(execute_CsrPlugin_csr_3008), .A2(
        _zz_CsrPlugin_csrMapping_readDataInit[28]), .B1(
        execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[28]), .ZN(n2255) );
  oai21d1 U3059 ( .B1(n3651), .B2(n2541), .A(n2255), .ZN(n2688) );
  inv0d0 U3060 ( .I(n2694), .ZN(n2683) );
  oai222d1 U3061 ( .A1(n2694), .A2(n2266), .B1(n2694), .B2(n2688), .C1(n2683), 
        .C2(n2289), .ZN(n3652) );
  oai22d1 U3062 ( .A1(n2256), .A2(n2303), .B1(n3652), .B2(n2322), .ZN(n6161)
         );
  inv0d0 U3063 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[27]), .ZN(n2258) );
  inv0d0 U3064 ( .I(CsrPlugin_mepc[27]), .ZN(n3648) );
  aoi22d1 U3065 ( .A1(execute_CsrPlugin_csr_3008), .A2(
        _zz_CsrPlugin_csrMapping_readDataInit[27]), .B1(
        execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[27]), .ZN(n2257) );
  oai21d1 U3066 ( .B1(n3648), .B2(n2541), .A(n2257), .ZN(n2693) );
  inv0d0 U3067 ( .I(n2711), .ZN(n2697) );
  oai222d1 U3068 ( .A1(n2711), .A2(n2266), .B1(n2711), .B2(n2693), .C1(n2697), 
        .C2(n2289), .ZN(n3649) );
  oai22d1 U3069 ( .A1(n2258), .A2(n2303), .B1(n3649), .B2(n2322), .ZN(n6160)
         );
  inv0d0 U3070 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[26]), .ZN(n2260) );
  aoi222d1 U3071 ( .A1(CsrPlugin_mepc[26]), .A2(execute_CsrPlugin_csr_833), 
        .B1(n2328), .B2(_zz_CsrPlugin_csrMapping_readDataInit[26]), .C1(n2327), 
        .C2(CsrPlugin_mtval[26]), .ZN(n2719) );
  inv0d0 U3072 ( .I(n2719), .ZN(n2259) );
  inv0d0 U3073 ( .I(n2713), .ZN(n2724) );
  oai222d1 U3074 ( .A1(n2713), .A2(n2266), .B1(n2713), .B2(n2259), .C1(n2724), 
        .C2(n2289), .ZN(n3646) );
  oai22d1 U3075 ( .A1(n2260), .A2(n2334), .B1(n3646), .B2(n2332), .ZN(n6159)
         );
  inv0d0 U3076 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[25]), .ZN(n2262) );
  aoi222d1 U3077 ( .A1(CsrPlugin_mepc[25]), .A2(execute_CsrPlugin_csr_833), 
        .B1(n2328), .B2(_zz_CsrPlugin_csrMapping_readDataInit[25]), .C1(n2327), 
        .C2(CsrPlugin_mtval[25]), .ZN(n2733) );
  inv0d0 U3078 ( .I(n2733), .ZN(n2261) );
  inv0d0 U3079 ( .I(n2728), .ZN(n2739) );
  oai222d1 U3080 ( .A1(n2728), .A2(n2266), .B1(n2728), .B2(n2261), .C1(n2739), 
        .C2(n2289), .ZN(n3643) );
  oai22d1 U3081 ( .A1(n2262), .A2(n2303), .B1(n3643), .B2(n2322), .ZN(n6158)
         );
  aoi222d1 U3082 ( .A1(CsrPlugin_mepc[24]), .A2(execute_CsrPlugin_csr_833), 
        .B1(n2328), .B2(_zz_CsrPlugin_csrMapping_readDataInit[24]), .C1(n2327), 
        .C2(CsrPlugin_mtval[24]), .ZN(n2747) );
  inv0d0 U3083 ( .I(n2747), .ZN(n2263) );
  inv0d0 U3084 ( .I(n2740), .ZN(n2754) );
  oai222d1 U3085 ( .A1(n2740), .A2(n2266), .B1(n2740), .B2(n2263), .C1(n2754), 
        .C2(n2331), .ZN(n3638) );
  inv0d0 U3086 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[24]), .ZN(n2264) );
  oai22d1 U3087 ( .A1(n3638), .A2(n2332), .B1(n2264), .B2(n2303), .ZN(n6157)
         );
  inv0d0 U3088 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[23]), .ZN(n2267) );
  inv0d0 U3089 ( .I(CsrPlugin_mepc[23]), .ZN(n3635) );
  aoi22d1 U3090 ( .A1(n2328), .A2(_zz_CsrPlugin_csrMapping_readDataInit[23]), 
        .B1(execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[23]), .ZN(n2265)
         );
  oai21d1 U3091 ( .B1(n3635), .B2(n2541), .A(n2265), .ZN(n2751) );
  inv0d0 U3092 ( .I(n2760), .ZN(n2755) );
  oai222d1 U3093 ( .A1(n2760), .A2(n2266), .B1(n2760), .B2(n2751), .C1(n2755), 
        .C2(n2289), .ZN(n3636) );
  oai22d1 U3094 ( .A1(n2267), .A2(n2334), .B1(n3636), .B2(n2332), .ZN(n6156)
         );
  aoi21d1 U3095 ( .B1(n2289), .B2(n2775), .A(n2269), .ZN(n3632) );
  inv0d0 U3096 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[22]), .ZN(n2270) );
  oai22d1 U3097 ( .A1(n3632), .A2(n2332), .B1(n2270), .B2(n2303), .ZN(n6155)
         );
  inv0d0 U3098 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[21]), .ZN(n2272) );
  inv0d0 U3099 ( .I(CsrPlugin_mepc[21]), .ZN(n3629) );
  aoi22d1 U3100 ( .A1(n2328), .A2(_zz_CsrPlugin_csrMapping_readDataInit[21]), 
        .B1(execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[21]), .ZN(n2271)
         );
  oai21d1 U3101 ( .B1(n3629), .B2(n2541), .A(n2271), .ZN(n2770) );
  inv0d0 U3102 ( .I(n2782), .ZN(n2790) );
  oai222d1 U3103 ( .A1(n2782), .A2(
        _zz__zz_execute_BranchPlugin_branch_src2[12]), .B1(n2782), .B2(n2770), 
        .C1(n2790), .C2(n2331), .ZN(n3630) );
  oai22d1 U3104 ( .A1(n2272), .A2(n2303), .B1(n3630), .B2(n2332), .ZN(n6154)
         );
  inv0d0 U3105 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[20]), .ZN(n2274) );
  inv0d0 U3106 ( .I(CsrPlugin_mepc[20]), .ZN(n3626) );
  aoi22d1 U3107 ( .A1(n2328), .A2(_zz_CsrPlugin_csrMapping_readDataInit[20]), 
        .B1(n2327), .B2(CsrPlugin_mtval[20]), .ZN(n2273) );
  oai21d1 U3108 ( .B1(n3626), .B2(n2541), .A(n2273), .ZN(n2785) );
  inv0d0 U3109 ( .I(n2805), .ZN(n2786) );
  oai222d1 U3110 ( .A1(n2805), .A2(n2266), .B1(n2805), .B2(n2785), .C1(n2786), 
        .C2(n2289), .ZN(n3627) );
  oai22d1 U3111 ( .A1(n2274), .A2(n2303), .B1(n3627), .B2(n2322), .ZN(n6153)
         );
  inv0d0 U3112 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[19]), .ZN(n2276) );
  inv0d0 U3113 ( .I(CsrPlugin_mepc[19]), .ZN(n3623) );
  aoi22d1 U3114 ( .A1(execute_CsrPlugin_csr_3008), .A2(
        _zz_CsrPlugin_csrMapping_readDataInit[19]), .B1(
        execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[19]), .ZN(n2275) );
  oai21d1 U3115 ( .B1(n3623), .B2(n2541), .A(n2275), .ZN(n2800) );
  inv0d0 U3116 ( .I(n2812), .ZN(n2819) );
  oai222d1 U3117 ( .A1(n2812), .A2(n2266), .B1(n2812), .B2(n2800), .C1(n2819), 
        .C2(n2331), .ZN(n3624) );
  oai22d1 U3118 ( .A1(n2276), .A2(n2334), .B1(n3624), .B2(n2322), .ZN(n6152)
         );
  inv0d0 U3119 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[18]), .ZN(n2278) );
  inv0d0 U3120 ( .I(CsrPlugin_mepc[18]), .ZN(n3620) );
  aoi22d1 U3121 ( .A1(n2328), .A2(_zz_CsrPlugin_csrMapping_readDataInit[18]), 
        .B1(execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[18]), .ZN(n2277)
         );
  oai21d1 U3122 ( .B1(n3620), .B2(n2541), .A(n2277), .ZN(n2823) );
  inv0d0 U3123 ( .I(n2835), .ZN(n2822) );
  oai222d1 U3124 ( .A1(n2835), .A2(n2266), .B1(n2835), .B2(n2823), .C1(n2822), 
        .C2(n2331), .ZN(n3621) );
  oai22d1 U3125 ( .A1(n2278), .A2(n2303), .B1(n3621), .B2(n2322), .ZN(n6151)
         );
  inv0d0 U3126 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[17]), .ZN(n2280) );
  inv0d0 U3127 ( .I(CsrPlugin_mepc[17]), .ZN(n3617) );
  aoi22d1 U3128 ( .A1(execute_CsrPlugin_csr_3008), .A2(
        _zz_CsrPlugin_csrMapping_readDataInit[17]), .B1(
        execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[17]), .ZN(n2279) );
  oai21d1 U3129 ( .B1(n3617), .B2(n2541), .A(n2279), .ZN(n2837) );
  inv0d0 U3130 ( .I(n2838), .ZN(n2836) );
  oai222d1 U3131 ( .A1(n2838), .A2(n2266), .B1(n2838), .B2(n2837), .C1(n2331), 
        .C2(n2836), .ZN(n3618) );
  oai22d1 U3132 ( .A1(n2280), .A2(n2303), .B1(n3618), .B2(n2332), .ZN(n6150)
         );
  inv0d0 U3133 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[16]), .ZN(n2283) );
  oai222d1 U3134 ( .A1(n2282), .A2(n2266), .B1(n2282), .B2(n2281), .C1(n2842), 
        .C2(n2289), .ZN(n3615) );
  oai22d1 U3135 ( .A1(n2283), .A2(n2334), .B1(n3615), .B2(n2332), .ZN(n6149)
         );
  inv0d0 U3136 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[15]), .ZN(n2286) );
  oai222d1 U3137 ( .A1(n2848), .A2(
        _zz__zz_execute_BranchPlugin_branch_src2[12]), .B1(n2848), .B2(n2285), 
        .C1(n2284), .C2(n2289), .ZN(n3612) );
  oai22d1 U3138 ( .A1(n2286), .A2(n2334), .B1(n3612), .B2(n2322), .ZN(n6148)
         );
  inv0d0 U3139 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[14]), .ZN(n2288) );
  inv0d0 U3140 ( .I(CsrPlugin_mepc[14]), .ZN(n3608) );
  aoi22d1 U3141 ( .A1(n2328), .A2(_zz_CsrPlugin_csrMapping_readDataInit[14]), 
        .B1(execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[14]), .ZN(n2287)
         );
  oai21d1 U3142 ( .B1(n3608), .B2(n2541), .A(n2287), .ZN(n2847) );
  oai222d1 U3143 ( .A1(n2863), .A2(n2266), .B1(n2863), .B2(n2847), .C1(n2860), 
        .C2(n2289), .ZN(n3609) );
  oai22d1 U3144 ( .A1(n2288), .A2(n2303), .B1(n3609), .B2(n2322), .ZN(n6147)
         );
  inv0d0 U3145 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[13]), .ZN(n2292) );
  oai222d1 U3146 ( .A1(n2291), .A2(
        _zz__zz_execute_BranchPlugin_branch_src2[12]), .B1(n2291), .B2(n2290), 
        .C1(n2855), .C2(n2289), .ZN(n3606) );
  oai22d1 U3147 ( .A1(n2292), .A2(n2303), .B1(n3606), .B2(n2322), .ZN(n6146)
         );
  inv0d0 U3148 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[12]), .ZN(n2295) );
  inv0d0 U3149 ( .I(n6919), .ZN(n2320) );
  oai222d1 U3150 ( .A1(n2869), .A2(n2320), .B1(n2869), .B2(n2294), .C1(n2293), 
        .C2(n2331), .ZN(n3603) );
  oai22d1 U3151 ( .A1(n2295), .A2(n2303), .B1(n3603), .B2(n2322), .ZN(n6145)
         );
  inv0d0 U3152 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[11]), .ZN(n2299) );
  aoi22d1 U3153 ( .A1(CsrPlugin_mepc[11]), .A2(execute_CsrPlugin_csr_833), 
        .B1(CsrPlugin_mstatus_MPP[0]), .B2(execute_CsrPlugin_csr_768), .ZN(
        n2298) );
  aoi22d1 U3154 ( .A1(execute_CsrPlugin_csr_3008), .A2(
        _zz_CsrPlugin_csrMapping_readDataInit[11]), .B1(CsrPlugin_mie_MEIE), 
        .B2(execute_CsrPlugin_csr_772), .ZN(n2297) );
  aoi22d1 U3155 ( .A1(n2327), .A2(CsrPlugin_mtval[11]), .B1(CsrPlugin_mip_MEIP), .B2(execute_CsrPlugin_csr_836), .ZN(n2296) );
  inv0d0 U3156 ( .I(n2873), .ZN(n2886) );
  oai222d1 U3157 ( .A1(n2873), .A2(n2320), .B1(n2873), .B2(n2871), .C1(n2331), 
        .C2(n2886), .ZN(n3600) );
  oai22d1 U3158 ( .A1(n2299), .A2(n2303), .B1(n3600), .B2(n2322), .ZN(n6144)
         );
  inv0d0 U3159 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[10]), .ZN(n2301) );
  inv0d0 U3160 ( .I(CsrPlugin_mepc[10]), .ZN(n3596) );
  aoi22d1 U3161 ( .A1(execute_CsrPlugin_csr_3008), .A2(
        _zz_CsrPlugin_csrMapping_readDataInit[10]), .B1(
        execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[10]), .ZN(n2300) );
  oai21d1 U3162 ( .B1(n3596), .B2(n2541), .A(n2300), .ZN(n2881) );
  inv0d0 U3163 ( .I(n2885), .ZN(n2900) );
  oai222d1 U3164 ( .A1(n2885), .A2(n2320), .B1(n2885), .B2(n2881), .C1(n2331), 
        .C2(n2900), .ZN(n3597) );
  oai22d1 U3165 ( .A1(n2301), .A2(n2334), .B1(n3597), .B2(n2322), .ZN(n6143)
         );
  inv0d0 U3166 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[9]), .ZN(n2304) );
  inv0d0 U3167 ( .I(CsrPlugin_mepc[9]), .ZN(n3593) );
  aoi22d1 U3168 ( .A1(execute_CsrPlugin_csr_3008), .A2(
        _zz_CsrPlugin_csrMapping_readDataInit[9]), .B1(
        execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[9]), .ZN(n2302) );
  oai21d1 U3169 ( .B1(n3593), .B2(n2541), .A(n2302), .ZN(n2904) );
  inv0d0 U3170 ( .I(n2899), .ZN(n2916) );
  oai222d1 U3171 ( .A1(n2899), .A2(n2320), .B1(n2899), .B2(n2904), .C1(n2331), 
        .C2(n2916), .ZN(n3594) );
  oai22d1 U3172 ( .A1(n2304), .A2(n2303), .B1(n3594), .B2(n2322), .ZN(n6142)
         );
  inv0d0 U3173 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[8]), .ZN(n2306) );
  inv0d0 U3174 ( .I(CsrPlugin_mepc[8]), .ZN(n3590) );
  aoi22d1 U3175 ( .A1(execute_CsrPlugin_csr_3008), .A2(
        _zz_CsrPlugin_csrMapping_readDataInit[8]), .B1(
        execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[8]), .ZN(n2305) );
  oai21d1 U3176 ( .B1(n3590), .B2(n2541), .A(n2305), .ZN(n2910) );
  inv0d0 U3177 ( .I(n2914), .ZN(n2933) );
  oai222d1 U3178 ( .A1(n2914), .A2(n2320), .B1(n2914), .B2(n2910), .C1(n2331), 
        .C2(n2933), .ZN(n3591) );
  oai22d1 U3179 ( .A1(n2306), .A2(n2334), .B1(n3591), .B2(n2322), .ZN(n6141)
         );
  inv0d0 U3180 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[7]), .ZN(n2311) );
  aoi22d1 U3181 ( .A1(CsrPlugin_mepc[7]), .A2(execute_CsrPlugin_csr_833), .B1(
        n2328), .B2(_zz_CsrPlugin_csrMapping_readDataInit[7]), .ZN(n2310) );
  aoi22d1 U3182 ( .A1(n2327), .A2(CsrPlugin_mtval[7]), .B1(
        execute_CsrPlugin_csr_768), .B2(CsrPlugin_mstatus_MPIE), .ZN(n2309) );
  aoi22d1 U3183 ( .A1(execute_CsrPlugin_csr_772), .A2(CsrPlugin_mie_MTIE), 
        .B1(n2307), .B2(execute_CsrPlugin_csr_4032), .ZN(n2308) );
  inv0d0 U3184 ( .I(n2931), .ZN(n2952) );
  oai222d1 U3185 ( .A1(n2931), .A2(n2320), .B1(n2931), .B2(n2926), .C1(n2331), 
        .C2(n2952), .ZN(n3588) );
  oai22d1 U3186 ( .A1(n2311), .A2(n2334), .B1(n3588), .B2(n2332), .ZN(n6140)
         );
  inv0d0 U3187 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[6]), .ZN(n2314) );
  aon211d1 U3188 ( .C1(execute_CsrPlugin_csr_4032), .C2(
        externalInterruptArray_regNext[6]), .B(execute_CsrPlugin_csr_3008), 
        .A(_zz_CsrPlugin_csrMapping_readDataInit[6]), .ZN(n2313) );
  aoi22d1 U3189 ( .A1(CsrPlugin_mepc[6]), .A2(execute_CsrPlugin_csr_833), .B1(
        execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[6]), .ZN(n2312) );
  nd02d0 U3190 ( .A1(n2313), .A2(n2312), .ZN(n2955) );
  inv0d0 U3191 ( .I(n2951), .ZN(n2966) );
  oai222d1 U3192 ( .A1(n2951), .A2(n2320), .B1(n2951), .B2(n2955), .C1(n2331), 
        .C2(n2966), .ZN(n3585) );
  oai22d1 U3193 ( .A1(n2314), .A2(n2334), .B1(n3585), .B2(n2332), .ZN(n6139)
         );
  inv0d0 U3194 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[5]), .ZN(n2317) );
  aoi22d1 U3195 ( .A1(CsrPlugin_mepc[5]), .A2(execute_CsrPlugin_csr_833), .B1(
        execute_CsrPlugin_csr_835), .B2(CsrPlugin_mtval[5]), .ZN(n2316) );
  aon211d1 U3196 ( .C1(execute_CsrPlugin_csr_4032), .C2(
        externalInterruptArray_regNext[5]), .B(execute_CsrPlugin_csr_3008), 
        .A(_zz_CsrPlugin_csrMapping_readDataInit[5]), .ZN(n2315) );
  nd02d0 U3197 ( .A1(n2316), .A2(n2315), .ZN(n2959) );
  inv0d0 U3198 ( .I(n2965), .ZN(n2981) );
  oai222d1 U3199 ( .A1(n2965), .A2(n2320), .B1(n2965), .B2(n2959), .C1(n2331), 
        .C2(n2981), .ZN(n3582) );
  oai22d1 U3200 ( .A1(n2317), .A2(n2334), .B1(n3582), .B2(n2332), .ZN(n6138)
         );
  inv0d0 U3201 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[4]), .ZN(n2321) );
  aoi22d1 U3202 ( .A1(CsrPlugin_mepc[4]), .A2(execute_CsrPlugin_csr_833), .B1(
        n2327), .B2(CsrPlugin_mtval[4]), .ZN(n2319) );
  aon211d1 U3203 ( .C1(execute_CsrPlugin_csr_4032), .C2(
        externalInterruptArray_regNext[4]), .B(execute_CsrPlugin_csr_3008), 
        .A(_zz_CsrPlugin_csrMapping_readDataInit[4]), .ZN(n2318) );
  nd02d0 U3204 ( .A1(n2319), .A2(n2318), .ZN(n2987) );
  oai222d1 U3205 ( .A1(n2990), .A2(n2320), .B1(n2990), .B2(n2987), .C1(n2985), 
        .C2(n2331), .ZN(n3579) );
  oai22d1 U3206 ( .A1(n2321), .A2(n2334), .B1(n3579), .B2(n2332), .ZN(n6137)
         );
  inv0d0 U3207 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[3]), .ZN(n2323) );
  inv0d0 U3208 ( .I(n2349), .ZN(n3576) );
  oai22d1 U3209 ( .A1(n2323), .A2(n2334), .B1(n3576), .B2(n2322), .ZN(n6136)
         );
  inv0d0 U3210 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[2]), .ZN(n2326) );
  inv0d0 U3211 ( .I(CsrPlugin_mtval[2]), .ZN(n2535) );
  aoi22d1 U3212 ( .A1(CsrPlugin_mepc[2]), .A2(execute_CsrPlugin_csr_833), .B1(
        execute_CsrPlugin_csr_834), .B2(CsrPlugin_mcause_exceptionCode[2]), 
        .ZN(n2325) );
  aon211d1 U3213 ( .C1(execute_CsrPlugin_csr_4032), .C2(
        externalInterruptArray_regNext[2]), .B(execute_CsrPlugin_csr_3008), 
        .A(_zz_CsrPlugin_csrMapping_readDataInit[2]), .ZN(n2324) );
  oai211d1 U3214 ( .C1(n2538), .C2(n2535), .A(n2325), .B(n2324), .ZN(n2998) );
  oai222d1 U3215 ( .A1(n3016), .A2(
        _zz__zz_execute_BranchPlugin_branch_src2[12]), .B1(n3016), .B2(n2998), 
        .C1(n2331), .C2(n3023), .ZN(n3573) );
  oai22d1 U3216 ( .A1(n2326), .A2(n2334), .B1(n3573), .B2(n2332), .ZN(n6135)
         );
  inv0d0 U3217 ( .I(_zz_CsrPlugin_csrMapping_readDataInit[1]), .ZN(n2333) );
  inv0d0 U3218 ( .I(CsrPlugin_mepc[1]), .ZN(n3569) );
  aoi22d1 U3219 ( .A1(execute_CsrPlugin_csr_834), .A2(
        CsrPlugin_mcause_exceptionCode[1]), .B1(n2327), .B2(CsrPlugin_mtval[1]), .ZN(n2330) );
  aon211d1 U3220 ( .C1(execute_CsrPlugin_csr_4032), .C2(
        externalInterruptArray_regNext[1]), .B(n2328), .A(
        _zz_CsrPlugin_csrMapping_readDataInit[1]), .ZN(n2329) );
  oai211d1 U3221 ( .C1(n2541), .C2(n3569), .A(n2330), .B(n2329), .ZN(n3021) );
  inv0d0 U3222 ( .I(n3039), .ZN(n3022) );
  oai222d1 U3223 ( .A1(n3039), .A2(
        _zz__zz_execute_BranchPlugin_branch_src2[12]), .B1(n3039), .B2(n3021), 
        .C1(n3022), .C2(n2331), .ZN(n3570) );
  oai22d1 U3224 ( .A1(n2334), .A2(n2333), .B1(n2332), .B2(n3570), .ZN(n6134)
         );
  aoim21d1 U3225 ( .B1(n2589), .B2(CsrPlugin_pipelineLiberator_pcValids_0), 
        .A(n2335), .ZN(n6131) );
  inv0d0 U3226 ( .I(CsrPlugin_mie_MEIE), .ZN(n2336) );
  inv0d0 U3227 ( .I(execute_CsrPlugin_csr_772), .ZN(n2545) );
  oai21d1 U3228 ( .B1(n3561), .B2(n2545), .A(n7121), .ZN(n2339) );
  nd03d0 U3229 ( .A1(n3566), .A2(execute_CsrPlugin_csr_772), .A3(n7121), .ZN(
        n2338) );
  oai22d1 U3230 ( .A1(n2336), .A2(n2339), .B1(n3600), .B2(n2338), .ZN(n6130)
         );
  inv0d0 U3231 ( .I(CsrPlugin_mie_MSIE), .ZN(n2337) );
  oai22d1 U3232 ( .A1(n2337), .A2(n2339), .B1(n3576), .B2(n2338), .ZN(n6129)
         );
  inv0d0 U3233 ( .I(CsrPlugin_mie_MTIE), .ZN(n2340) );
  oai22d1 U3234 ( .A1(n2340), .A2(n2339), .B1(n3588), .B2(n2338), .ZN(n6128)
         );
  nd02d0 U3235 ( .A1(n3566), .A2(execute_CsrPlugin_csr_768), .ZN(n2348) );
  nd02d0 U3236 ( .A1(n2393), .A2(n2348), .ZN(n2345) );
  nd02d0 U3237 ( .A1(n7121), .A2(n2345), .ZN(n2353) );
  inv0d0 U3238 ( .I(n2353), .ZN(n2344) );
  inv0d0 U3239 ( .I(n2351), .ZN(n2342) );
  oan211d1 U3240 ( .C1(n2348), .C2(n3600), .B(n2344), .A(n2341), .ZN(n6127) );
  nr02d0 U3241 ( .A1(CsrPlugin_mstatus_MPP[1]), .A2(n2342), .ZN(n2343) );
  oan211d1 U3242 ( .C1(n2348), .C2(n3603), .B(n2344), .A(n2343), .ZN(n6126) );
  inv0d0 U3243 ( .I(n2348), .ZN(n2350) );
  aon211d1 U3244 ( .C1(CsrPlugin_mstatus_MIE), .C2(n3672), .B(n2345), .A(n7121), .ZN(n2347) );
  nd02d0 U3245 ( .A1(n2351), .A2(CsrPlugin_mstatus_MPIE), .ZN(n2346) );
  aon211d1 U3246 ( .C1(n2350), .C2(n3588), .B(n2347), .A(n2346), .ZN(n6125) );
  aoi22d1 U3247 ( .A1(n2350), .A2(n2349), .B1(CsrPlugin_mstatus_MPIE), .B2(
        n2348), .ZN(n2352) );
  oaim22d1 U3248 ( .A1(n2353), .A2(n2352), .B1(n2351), .B2(
        CsrPlugin_mstatus_MIE), .ZN(n6124) );
  inv0d0 U3249 ( .I(n3697), .ZN(n3687) );
  nr02d0 U3250 ( .A1(n2354), .A2(n3687), .ZN(n3694) );
  aoi211d1 U3251 ( .C1(n3679), .C2(n3687), .A(n3694), .B(n2355), .ZN(n6123) );
  inv0d0 U3252 ( .I(n2356), .ZN(n6908) );
  inv0d2 U3253 ( .I(n6893), .ZN(n6862) );
  aoi221d1 U3254 ( .B1(n7007), .B2(n2372), .C1(n6862), .C2(n2359), .A(n2373), 
        .ZN(n6120) );
  aor31d1 U3255 ( .B1(n2361), .B2(n2360), .B3(n2577), .A(
        \IBusCachedPlugin_cache/lineLoader_flushPending ), .Z(n2411) );
  inv0d0 U3256 ( .I(n2362), .ZN(n2366) );
  nr02d0 U3257 ( .A1(n2412), .A2(n3287), .ZN(n2364) );
  inv0d0 U3258 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port[0] ), .ZN(
        n3054) );
  nr04d0 U3259 ( .A1(DebugPlugin_haltIt), .A2(CsrPlugin_exceptionPendings_3), 
        .A3(\IBusCachedPlugin_cache/lineLoader_valid ), .A4(n3054), .ZN(n2363)
         );
  oai21d1 U3260 ( .B1(IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid), 
        .B2(_zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1), .A(
        DebugPlugin_stepIt), .ZN(n2425) );
  nr04d0 U3261 ( .A1(n2367), .A2(n2411), .A3(n2366), .A4(n2365), .ZN(n2371) );
  inv0d0 U3262 ( .I(n2368), .ZN(n2370) );
  oai31d1 U3263 ( .B1(n3818), .B2(n2373), .B3(n2372), .A(n2375), .ZN(n6119) );
  nd02d0 U3264 ( .A1(n2397), .A2(n2374), .ZN(n2377) );
  inv0d0 U3265 ( .I(\_zz_IBusCachedPlugin_fetchPc_pc_1[2] ), .ZN(n2376) );
  oai31d1 U3266 ( .B1(reset), .B2(n2377), .B3(n2376), .A(n2375), .ZN(n6118) );
  aoi22d1 U3267 ( .A1(n2394), .A2(CsrPlugin_mepc[2]), .B1(
        CsrPlugin_mtvec_base[0]), .B2(n2393), .ZN(n2381) );
  ah01d1 U3268 ( .A(IBusCachedPlugin_iBusRsp_stages_1_input_payload[2]), .B(
        \_zz_IBusCachedPlugin_fetchPc_pc_1[2] ), .CO(n2383), .S(n2378) );
  aoi22d1 U3269 ( .A1(n2398), .A2(memory_BRANCH_CALC[2]), .B1(n2397), .B2(
        n2378), .ZN(n2380) );
  nd02d0 U3270 ( .A1(n2399), .A2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[2]), .ZN(
        n2379) );
  oai211d1 U3271 ( .C1(n2403), .C2(n2381), .A(n2380), .B(n2379), .ZN(n3706) );
  inv0d0 U3272 ( .I(n3706), .ZN(n3709) );
  inv0d0 U3273 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[2]), .ZN(
        n3246) );
  inv0d0 U3274 ( .I(n2382), .ZN(n2404) );
  oai22d1 U3275 ( .A1(n3709), .A2(n2405), .B1(n3246), .B2(n2404), .ZN(n6117)
         );
  aoi22d1 U3276 ( .A1(n2394), .A2(CsrPlugin_mepc[3]), .B1(
        CsrPlugin_mtvec_base[1]), .B2(n2393), .ZN(n2386) );
  ah01d1 U3277 ( .A(n2383), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[3]), .CO(n2388), .S(
        n2384) );
  aoi22d1 U3278 ( .A1(n2398), .A2(memory_BRANCH_CALC[3]), .B1(n2397), .B2(
        n2384), .ZN(n2385) );
  oai21d1 U3279 ( .B1(n2403), .B2(n2386), .A(n2385), .ZN(n2387) );
  aoi21d1 U3280 ( .B1(n2399), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[3]), .A(n2387), .ZN(n3705) );
  inv0d0 U3281 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[3]), .ZN(
        n3242) );
  oai22d1 U3282 ( .A1(n3705), .A2(n2405), .B1(n3242), .B2(n2404), .ZN(n6116)
         );
  aoi22d1 U3283 ( .A1(n2394), .A2(CsrPlugin_mepc[4]), .B1(
        CsrPlugin_mtvec_base[2]), .B2(n2393), .ZN(n2391) );
  ah01d1 U3284 ( .A(n2388), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[4]), .CO(n2395), .S(
        n2389) );
  aoi22d1 U3285 ( .A1(n2399), .A2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[4]), .B1(
        n2397), .B2(n2389), .ZN(n2390) );
  oai21d1 U3286 ( .B1(n2403), .B2(n2391), .A(n2390), .ZN(n2392) );
  aoi21d1 U3287 ( .B1(n2398), .B2(memory_BRANCH_CALC[4]), .A(n2392), .ZN(n3710) );
  inv0d0 U3288 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[4]), .ZN(
        n3240) );
  oai22d1 U3289 ( .A1(n3710), .A2(n2405), .B1(n3240), .B2(n2404), .ZN(n6115)
         );
  aoi22d1 U3290 ( .A1(n2394), .A2(CsrPlugin_mepc[5]), .B1(
        CsrPlugin_mtvec_base[3]), .B2(n2393), .ZN(n2402) );
  ah01d1 U3291 ( .A(n2395), .B(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[5]), .CO(n452), .S(
        n2396) );
  aoi22d1 U3292 ( .A1(n2398), .A2(memory_BRANCH_CALC[5]), .B1(n2397), .B2(
        n2396), .ZN(n2401) );
  nd02d0 U3293 ( .A1(n2399), .A2(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[5]), .ZN(
        n2400) );
  oai211d1 U3294 ( .C1(n2403), .C2(n2402), .A(n2401), .B(n2400), .ZN(n7005) );
  inv0d0 U3295 ( .I(n7005), .ZN(n7006) );
  inv0d0 U3296 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[5]), .ZN(
        n7001) );
  oai22d1 U3297 ( .A1(n7006), .A2(n2405), .B1(n7001), .B2(n2404), .ZN(n6114)
         );
  aon211d1 U3298 ( .C1(\IBusCachedPlugin_cache/lineLoader_flushCounter[0] ), 
        .C2(\IBusCachedPlugin_cache/_zz_ways_0_tags_port[0] ), .B(n3060), .A(
        n2410), .ZN(n2406) );
  inv0d0 U3299 ( .I(n2406), .ZN(n6087) );
  inv0d0 U3300 ( .I(n2407), .ZN(n3059) );
  aoim211d1 U3301 ( .C1(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[0] ), 
        .C2(iBus_rsp_valid), .A(reset), .B(n3059), .ZN(n6085) );
  inv0d0 U3302 ( .I(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[1] ), 
        .ZN(n3159) );
  aoi221d1 U3303 ( .B1(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[1] ), 
        .B2(n3059), .C1(n3159), .C2(n2407), .A(reset), .ZN(n6084) );
  inv0d0 U3304 ( .I(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[2] ), 
        .ZN(n2409) );
  nd02d0 U3305 ( .A1(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[1] ), 
        .A2(n3059), .ZN(n2408) );
  aoi211d1 U3306 ( .C1(n2409), .C2(n2408), .A(reset), .B(n2414), .ZN(n6083) );
  oaim21d1 U3307 ( .B1(n2411), .B2(n2410), .A(n7121), .ZN(n6081) );
  oan211d1 U3308 ( .C1(n2414), .C2(n2413), .B(n3049), .A(n2412), .ZN(n6080) );
  nd12d0 U3309 ( .A1(debug_bus_cmd_payload_address[2]), .A2(n2415), .ZN(n2423)
         );
  inv0d0 U3310 ( .I(n2423), .ZN(n3703) );
  inv0d0 U3311 ( .I(debugReset), .ZN(n3701) );
  aon211d1 U3312 ( .C1(debug_bus_cmd_payload_data[18]), .C2(n3703), .B(
        DebugPlugin_disableEbreak), .A(n3701), .ZN(n2416) );
  aoi21d1 U3313 ( .B1(debug_bus_cmd_payload_data[26]), .B2(n3703), .A(n2416), 
        .ZN(n6079) );
  aoim21d1 U3314 ( .B1(debug_bus_cmd_valid), .B2(DebugPlugin_debugUsed), .A(
        debugReset), .ZN(n6078) );
  nr02d0 U3315 ( .A1(n2420), .A2(n2423), .ZN(n2419) );
  nd02d0 U3316 ( .A1(n2428), .A2(n2427), .ZN(n2417) );
  oan211d1 U3317 ( .C1(n2419), .C2(n2418), .B(n2417), .A(debugReset), .ZN(
        n6077) );
  inv0d0 U3318 ( .I(DebugPlugin_godmode), .ZN(n2421) );
  oai21d1 U3319 ( .B1(n2420), .B2(n2423), .A(n3701), .ZN(n2430) );
  oan211d1 U3320 ( .C1(DebugPlugin_isPipBusy), .C2(n2435), .B(n2421), .A(n2430), .ZN(n6076) );
  aoi221d1 U3321 ( .B1(n3703), .B2(n2424), .C1(n2423), .C2(n2422), .A(
        debugReset), .ZN(n6075) );
  aoim22d1 U3322 ( .A1(n2428), .A2(n2427), .B1(n2426), .B2(n2425), .Z(n2429)
         );
  inv0d0 U3323 ( .I(n2429), .ZN(n2431) );
  aoi211d1 U3324 ( .C1(debug_bus_cmd_payload_data[17]), .C2(n3703), .A(n2431), 
        .B(n2430), .ZN(n2432) );
  mx02d1 U3325 ( .I0(n2433), .I1(DebugPlugin_haltIt), .S(n2432), .Z(n6074) );
  nd03d0 U3326 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[6]), .A2(
        _zz_decode_LEGAL_INSTRUCTION_1[4]), .A3(n2434), .ZN(n2560) );
  nr03d0 U3327 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13[28]), .A2(n3238), .A3(
        n2560), .ZN(n2562) );
  nd04d0 U3328 ( .A1(\_zz__zz_decode_ENV_CTRL_2_1[20] ), .A2(n2562), .A3(
        DebugPlugin_debugUsed), .A4(n2435), .ZN(n2436) );
  oaim22d1 U3329 ( .A1(DebugPlugin_disableEbreak), .A2(n2436), .B1(n3235), 
        .B2(execute_DO_EBREAK), .ZN(n6073) );
  aoi22d1 U3330 ( .A1(n2483), .A2(iBus_rsp_payload_data[18]), .B1(n2458), .B2(
        iBus_rsp_payload_data[10]), .ZN(n2439) );
  aoi22d1 U3331 ( .A1(n2462), .A2(iBus_rsp_payload_data[2]), .B1(n2453), .B2(
        iBus_rsp_payload_data[26]), .ZN(n2438) );
  nd02d0 U3332 ( .A1(n2526), .A2(writeBack_REGFILE_WRITE_DATA[2]), .ZN(n2437)
         );
  aon211d1 U3333 ( .C1(n2439), .C2(n2438), .B(n2526), .A(n2437), .ZN(n3284) );
  inv0d0 U3334 ( .I(n3284), .ZN(n3427) );
  inv0d0 U3335 ( .I(execute_PC[2]), .ZN(n6299) );
  oai222d1 U3336 ( .A1(n2440), .A2(n2514), .B1(n2531), .B2(n3427), .C1(n2530), 
        .C2(n6299), .ZN(n6070) );
  aoi22d1 U3337 ( .A1(n2453), .A2(iBus_rsp_payload_data[27]), .B1(n2483), .B2(
        iBus_rsp_payload_data[19]), .ZN(n2443) );
  aoi22d1 U3338 ( .A1(n2462), .A2(iBus_rsp_payload_data[3]), .B1(n2458), .B2(
        iBus_rsp_payload_data[11]), .ZN(n2442) );
  nd02d0 U3339 ( .A1(n2526), .A2(writeBack_REGFILE_WRITE_DATA[3]), .ZN(n2441)
         );
  aon211d1 U3340 ( .C1(n2443), .C2(n2442), .B(n2526), .A(n2441), .ZN(n3283) );
  inv0d0 U3341 ( .I(n3283), .ZN(n3424) );
  inv0d0 U3342 ( .I(execute_PC[3]), .ZN(n6420) );
  oai222d1 U3343 ( .A1(n2444), .A2(n2514), .B1(n2531), .B2(n3424), .C1(n2530), 
        .C2(n6420), .ZN(n6069) );
  buffd1 U3344 ( .I(n2514), .Z(n2532) );
  aoi22d1 U3345 ( .A1(n2453), .A2(iBus_rsp_payload_data[28]), .B1(n2458), .B2(
        iBus_rsp_payload_data[12]), .ZN(n2447) );
  aoi22d1 U3346 ( .A1(n2462), .A2(iBus_rsp_payload_data[4]), .B1(n2483), .B2(
        iBus_rsp_payload_data[20]), .ZN(n2446) );
  nd02d0 U3347 ( .A1(n2526), .A2(writeBack_REGFILE_WRITE_DATA[4]), .ZN(n2445)
         );
  aon211d1 U3348 ( .C1(n2447), .C2(n2446), .B(n2526), .A(n2445), .ZN(n3281) );
  inv0d0 U3349 ( .I(n3281), .ZN(n3423) );
  inv0d0 U3350 ( .I(execute_PC[4]), .ZN(n7114) );
  oai222d1 U3351 ( .A1(n2448), .A2(n2532), .B1(n2531), .B2(n3423), .C1(n2530), 
        .C2(n7114), .ZN(n6068) );
  inv0d0 U3352 ( .I(debug_bus_rsp_data[5]), .ZN(n2452) );
  aoi22d1 U3353 ( .A1(n2462), .A2(iBus_rsp_payload_data[5]), .B1(n2483), .B2(
        iBus_rsp_payload_data[21]), .ZN(n2451) );
  aoi22d1 U3354 ( .A1(n2453), .A2(iBus_rsp_payload_data[29]), .B1(n2458), .B2(
        iBus_rsp_payload_data[13]), .ZN(n2450) );
  nd02d0 U3355 ( .A1(n2526), .A2(writeBack_REGFILE_WRITE_DATA[5]), .ZN(n2449)
         );
  aon211d1 U3356 ( .C1(n2451), .C2(n2450), .B(n2526), .A(n2449), .ZN(n3280) );
  inv0d0 U3357 ( .I(n3280), .ZN(n3422) );
  inv0d0 U3358 ( .I(execute_PC[5]), .ZN(n7002) );
  oai222d1 U3359 ( .A1(n2452), .A2(n2532), .B1(n2531), .B2(n3422), .C1(n2530), 
        .C2(n7002), .ZN(n6067) );
  inv0d0 U3360 ( .I(debug_bus_rsp_data[6]), .ZN(n2457) );
  aoi22d1 U3361 ( .A1(n2453), .A2(iBus_rsp_payload_data[30]), .B1(n2483), .B2(
        iBus_rsp_payload_data[22]), .ZN(n2456) );
  aoi22d1 U3362 ( .A1(n2462), .A2(iBus_rsp_payload_data[6]), .B1(n2458), .B2(
        iBus_rsp_payload_data[14]), .ZN(n2455) );
  nd02d0 U3363 ( .A1(n2526), .A2(writeBack_REGFILE_WRITE_DATA[6]), .ZN(n2454)
         );
  aon211d1 U3364 ( .C1(n2456), .C2(n2455), .B(n2526), .A(n2454), .ZN(n3278) );
  inv0d0 U3365 ( .I(n3278), .ZN(n3421) );
  inv0d0 U3366 ( .I(execute_PC[6]), .ZN(n6940) );
  oai222d1 U3367 ( .A1(n2457), .A2(n2514), .B1(n2531), .B2(n3421), .C1(n2474), 
        .C2(n6940), .ZN(n6066) );
  inv0d0 U3368 ( .I(debug_bus_rsp_data[7]), .ZN(n2463) );
  aoi22d1 U3369 ( .A1(n2483), .A2(iBus_rsp_payload_data[23]), .B1(n2458), .B2(
        iBus_rsp_payload_data[15]), .ZN(n2459) );
  oai21d1 U3370 ( .B1(n2460), .B2(n3166), .A(n2459), .ZN(n2461) );
  aon211d1 U3371 ( .C1(n2462), .C2(iBus_rsp_payload_data[7]), .B(n2461), .A(
        n2476), .ZN(n2464) );
  oaim21d1 U3372 ( .B1(writeBack_REGFILE_WRITE_DATA[7]), .B2(n2526), .A(n2464), 
        .ZN(n3277) );
  inv0d0 U3373 ( .I(n3277), .ZN(n3420) );
  inv0d0 U3374 ( .I(execute_PC[7]), .ZN(n6927) );
  oai222d1 U3375 ( .A1(n2463), .A2(n2514), .B1(n2531), .B2(n3420), .C1(n2474), 
        .C2(n6927), .ZN(n6065) );
  inv0d0 U3376 ( .I(debug_bus_rsp_data[8]), .ZN(n2466) );
  an02d0 U3377 ( .A1(n2476), .A2(_zz_lastStageRegFileWrite_payload_address[12]), .Z(n2491) );
  an02d1 U3378 ( .A1(n2476), .A2(_zz_lastStageRegFileWrite_payload_address[13]), .Z(n2527) );
  buffd1 U3379 ( .I(n2527), .Z(n2523) );
  oai21d1 U3380 ( .B1(n2491), .B2(n2523), .A(n2483), .ZN(n2481) );
  nr02d0 U3381 ( .A1(n2491), .A2(n2523), .ZN(n2484) );
  aoi22d1 U3382 ( .A1(iBus_rsp_payload_data[8]), .A2(n2479), .B1(
        writeBack_REGFILE_WRITE_DATA[8]), .B2(n2526), .ZN(n2465) );
  nr04d0 U3383 ( .A1(_zz_lastStageRegFileWrite_payload_address[14]), .A2(
        _zz_lastStageRegFileWrite_payload_address[12]), .A3(
        _zz_lastStageRegFileWrite_payload_address[13]), .A4(n2464), .ZN(n2489)
         );
  inv0d0 U3384 ( .I(n2489), .ZN(n2486) );
  oai211d1 U3385 ( .C1(n3179), .C2(n2481), .A(n2465), .B(n2486), .ZN(n3276) );
  inv0d0 U3386 ( .I(n3276), .ZN(n3419) );
  inv0d0 U3387 ( .I(execute_PC[8]), .ZN(n6916) );
  oai222d1 U3388 ( .A1(n2466), .A2(n2514), .B1(n2531), .B2(n3419), .C1(n2474), 
        .C2(n6916), .ZN(n6064) );
  inv0d0 U3389 ( .I(debug_bus_rsp_data[9]), .ZN(n2468) );
  aoi22d1 U3390 ( .A1(iBus_rsp_payload_data[9]), .A2(n2479), .B1(
        writeBack_REGFILE_WRITE_DATA[9]), .B2(n2526), .ZN(n2467) );
  oai211d1 U3391 ( .C1(n3178), .C2(n2481), .A(n2467), .B(n2486), .ZN(n3275) );
  inv0d0 U3392 ( .I(n3275), .ZN(n3418) );
  inv0d0 U3393 ( .I(execute_PC[9]), .ZN(n6911) );
  oai222d1 U3394 ( .A1(n2468), .A2(n2532), .B1(n2531), .B2(n3418), .C1(n2474), 
        .C2(n6911), .ZN(n6063) );
  inv0d0 U3395 ( .I(debug_bus_rsp_data[10]), .ZN(n2470) );
  aoi22d1 U3396 ( .A1(iBus_rsp_payload_data[10]), .A2(n2479), .B1(
        writeBack_REGFILE_WRITE_DATA[10]), .B2(n2526), .ZN(n2469) );
  oai211d1 U3397 ( .C1(n3177), .C2(n2481), .A(n2469), .B(n2486), .ZN(n3274) );
  inv0d0 U3398 ( .I(n3274), .ZN(n3417) );
  inv0d0 U3399 ( .I(execute_PC[10]), .ZN(n6905) );
  oai222d1 U3400 ( .A1(n2470), .A2(n2532), .B1(n2531), .B2(n3417), .C1(n2474), 
        .C2(n6905), .ZN(n6062) );
  inv0d0 U3401 ( .I(debug_bus_rsp_data[11]), .ZN(n2472) );
  aoi22d1 U3402 ( .A1(iBus_rsp_payload_data[11]), .A2(n2479), .B1(
        writeBack_REGFILE_WRITE_DATA[11]), .B2(n2526), .ZN(n2471) );
  oai211d1 U3403 ( .C1(n3176), .C2(n2481), .A(n2471), .B(n2486), .ZN(n3273) );
  inv0d0 U3404 ( .I(n3273), .ZN(n3416) );
  inv0d0 U3405 ( .I(execute_PC[11]), .ZN(n6900) );
  oai222d1 U3406 ( .A1(n2472), .A2(n2532), .B1(n2531), .B2(n3416), .C1(n2474), 
        .C2(n6900), .ZN(n6061) );
  inv0d0 U3407 ( .I(debug_bus_rsp_data[12]), .ZN(n2475) );
  aoi22d1 U3408 ( .A1(iBus_rsp_payload_data[12]), .A2(n2479), .B1(
        writeBack_REGFILE_WRITE_DATA[12]), .B2(n2526), .ZN(n2473) );
  oai211d1 U3409 ( .C1(n3175), .C2(n2481), .A(n2473), .B(n2486), .ZN(n3272) );
  inv0d0 U3410 ( .I(n3272), .ZN(n3415) );
  inv0d0 U3411 ( .I(execute_PC[12]), .ZN(n7118) );
  oai222d1 U3412 ( .A1(n2475), .A2(n2532), .B1(n2531), .B2(n3415), .C1(n2474), 
        .C2(n7118), .ZN(n6060) );
  inv0d0 U3413 ( .I(debug_bus_rsp_data[13]), .ZN(n2478) );
  inv0d1 U3414 ( .I(n2476), .ZN(n2522) );
  aoi22d1 U3415 ( .A1(iBus_rsp_payload_data[13]), .A2(n2479), .B1(
        writeBack_REGFILE_WRITE_DATA[13]), .B2(n2522), .ZN(n2477) );
  oai211d1 U3416 ( .C1(n3174), .C2(n2481), .A(n2477), .B(n2486), .ZN(n3271) );
  inv0d0 U3417 ( .I(n3271), .ZN(n3414) );
  inv0d0 U3418 ( .I(execute_PC[13]), .ZN(n6894) );
  oai222d1 U3419 ( .A1(n2478), .A2(n2532), .B1(n2531), .B2(n3414), .C1(n2530), 
        .C2(n6894), .ZN(n6059) );
  inv0d0 U3420 ( .I(debug_bus_rsp_data[14]), .ZN(n2482) );
  aoi22d1 U3421 ( .A1(n2479), .A2(iBus_rsp_payload_data[14]), .B1(
        writeBack_REGFILE_WRITE_DATA[14]), .B2(n2522), .ZN(n2480) );
  oai211d1 U3422 ( .C1(n3173), .C2(n2481), .A(n2480), .B(n2486), .ZN(n3270) );
  inv0d0 U3423 ( .I(n3270), .ZN(n3413) );
  inv0d0 U3424 ( .I(execute_PC[14]), .ZN(n6887) );
  oai222d1 U3425 ( .A1(n2482), .A2(n2514), .B1(n2531), .B2(n3413), .C1(n2530), 
        .C2(n6887), .ZN(n6058) );
  inv0d0 U3426 ( .I(debug_bus_rsp_data[15]), .ZN(n2488) );
  aoim22d1 U3427 ( .A1(n2483), .A2(n3166), .B1(iBus_rsp_payload_data[15]), 
        .B2(n2483), .Z(n2490) );
  inv0d0 U3428 ( .I(n2484), .ZN(n2485) );
  aoi22d1 U3429 ( .A1(writeBack_REGFILE_WRITE_DATA[15]), .A2(n2522), .B1(n2490), .B2(n2485), .ZN(n2487) );
  nd02d0 U3430 ( .A1(n2487), .A2(n2486), .ZN(n3269) );
  inv0d0 U3431 ( .I(n3269), .ZN(n3412) );
  inv0d0 U3432 ( .I(execute_PC[15]), .ZN(n6882) );
  oai222d1 U3433 ( .A1(n2488), .A2(n2514), .B1(n2531), .B2(n3412), .C1(n2530), 
        .C2(n6882), .ZN(n6057) );
  inv0d0 U3434 ( .I(debug_bus_rsp_data[16]), .ZN(n2494) );
  nr02d0 U3435 ( .A1(_zz_lastStageRegFileWrite_payload_address[14]), .A2(
        _zz_lastStageRegFileWrite_payload_address[13]), .ZN(n2492) );
  aoi31d1 U3436 ( .B1(n2492), .B2(n2491), .B3(n2490), .A(n2489), .ZN(n2529) );
  aoi22d1 U3437 ( .A1(iBus_rsp_payload_data[16]), .A2(n2527), .B1(
        writeBack_REGFILE_WRITE_DATA[16]), .B2(n2522), .ZN(n2493) );
  nd02d0 U3438 ( .A1(n2529), .A2(n2493), .ZN(n3268) );
  inv0d0 U3439 ( .I(n3268), .ZN(n3411) );
  inv0d0 U3440 ( .I(execute_PC[16]), .ZN(n6875) );
  oai222d1 U3441 ( .A1(n2494), .A2(n2532), .B1(n2531), .B2(n3411), .C1(n2530), 
        .C2(n6875), .ZN(n6056) );
  inv0d0 U3442 ( .I(debug_bus_rsp_data[17]), .ZN(n2496) );
  aoi22d1 U3443 ( .A1(iBus_rsp_payload_data[17]), .A2(n2527), .B1(
        writeBack_REGFILE_WRITE_DATA[17]), .B2(n2522), .ZN(n2495) );
  nd02d0 U3444 ( .A1(n2529), .A2(n2495), .ZN(n3267) );
  inv0d0 U3445 ( .I(n3267), .ZN(n3410) );
  inv0d0 U3446 ( .I(execute_PC[17]), .ZN(n6870) );
  oai222d1 U3447 ( .A1(n2496), .A2(n2514), .B1(n2531), .B2(n3410), .C1(n2530), 
        .C2(n6870), .ZN(n6055) );
  inv0d0 U3448 ( .I(debug_bus_rsp_data[18]), .ZN(n2498) );
  aoi22d1 U3449 ( .A1(iBus_rsp_payload_data[18]), .A2(n2527), .B1(
        writeBack_REGFILE_WRITE_DATA[18]), .B2(n2522), .ZN(n2497) );
  nd02d0 U3450 ( .A1(n2529), .A2(n2497), .ZN(n3266) );
  inv0d0 U3451 ( .I(n3266), .ZN(n3409) );
  inv0d0 U3452 ( .I(execute_PC[18]), .ZN(n6865) );
  oai222d1 U3453 ( .A1(n2498), .A2(n2514), .B1(n2531), .B2(n3409), .C1(n2530), 
        .C2(n6865), .ZN(n6054) );
  inv0d0 U3454 ( .I(debug_bus_rsp_data[19]), .ZN(n2500) );
  aoi22d1 U3455 ( .A1(iBus_rsp_payload_data[19]), .A2(n2527), .B1(
        writeBack_REGFILE_WRITE_DATA[19]), .B2(n2522), .ZN(n2499) );
  nd02d0 U3456 ( .A1(n2529), .A2(n2499), .ZN(n3265) );
  inv0d0 U3457 ( .I(n3265), .ZN(n3408) );
  inv0d0 U3458 ( .I(execute_PC[19]), .ZN(n6859) );
  oai222d1 U3459 ( .A1(n2500), .A2(n2532), .B1(n2531), .B2(n3408), .C1(n2530), 
        .C2(n6859), .ZN(n6053) );
  inv0d0 U3460 ( .I(debug_bus_rsp_data[20]), .ZN(n2502) );
  aoi22d1 U3461 ( .A1(iBus_rsp_payload_data[20]), .A2(n2527), .B1(
        writeBack_REGFILE_WRITE_DATA[20]), .B2(n2522), .ZN(n2501) );
  nd02d0 U3462 ( .A1(n2529), .A2(n2501), .ZN(n3264) );
  inv0d0 U3463 ( .I(n3264), .ZN(n3407) );
  inv0d0 U3464 ( .I(execute_PC[20]), .ZN(n6854) );
  oai222d1 U3465 ( .A1(n2502), .A2(n2514), .B1(n2531), .B2(n3407), .C1(n2530), 
        .C2(n6854), .ZN(n6052) );
  inv0d0 U3466 ( .I(debug_bus_rsp_data[21]), .ZN(n2504) );
  aoi22d1 U3467 ( .A1(iBus_rsp_payload_data[21]), .A2(n2527), .B1(
        writeBack_REGFILE_WRITE_DATA[21]), .B2(n2522), .ZN(n2503) );
  nd02d0 U3468 ( .A1(n2529), .A2(n2503), .ZN(n3263) );
  inv0d0 U3469 ( .I(n3263), .ZN(n3406) );
  inv0d0 U3470 ( .I(execute_PC[21]), .ZN(n6849) );
  oai222d1 U3471 ( .A1(n2504), .A2(n2532), .B1(n2531), .B2(n3406), .C1(n2530), 
        .C2(n6849), .ZN(n6051) );
  inv0d0 U3472 ( .I(debug_bus_rsp_data[22]), .ZN(n2506) );
  aoi22d1 U3473 ( .A1(iBus_rsp_payload_data[22]), .A2(n2527), .B1(
        writeBack_REGFILE_WRITE_DATA[22]), .B2(n2522), .ZN(n2505) );
  nd02d0 U3474 ( .A1(n2529), .A2(n2505), .ZN(n3262) );
  inv0d0 U3475 ( .I(n3262), .ZN(n3405) );
  inv0d0 U3476 ( .I(execute_PC[22]), .ZN(n6844) );
  oai222d1 U3477 ( .A1(n2506), .A2(n2514), .B1(n2531), .B2(n3405), .C1(n2530), 
        .C2(n6844), .ZN(n6050) );
  inv0d0 U3478 ( .I(debug_bus_rsp_data[23]), .ZN(n2508) );
  aoi22d1 U3479 ( .A1(n2527), .A2(iBus_rsp_payload_data[23]), .B1(
        writeBack_REGFILE_WRITE_DATA[23]), .B2(n2522), .ZN(n2507) );
  nd02d0 U3480 ( .A1(n2529), .A2(n2507), .ZN(n3261) );
  inv0d0 U3481 ( .I(n3261), .ZN(n3404) );
  inv0d0 U3482 ( .I(execute_PC[23]), .ZN(n6839) );
  oai222d1 U3483 ( .A1(n2508), .A2(n2532), .B1(n2531), .B2(n3404), .C1(n2530), 
        .C2(n6839), .ZN(n6049) );
  inv0d0 U3484 ( .I(debug_bus_rsp_data[24]), .ZN(n2510) );
  aoi22d1 U3485 ( .A1(iBus_rsp_payload_data[24]), .A2(n2523), .B1(
        writeBack_REGFILE_WRITE_DATA[24]), .B2(n2522), .ZN(n2509) );
  nd02d0 U3486 ( .A1(n2529), .A2(n2509), .ZN(n3260) );
  inv0d0 U3487 ( .I(n3260), .ZN(n3403) );
  inv0d0 U3488 ( .I(execute_PC[24]), .ZN(n6834) );
  oai222d1 U3489 ( .A1(n2510), .A2(n2532), .B1(n2531), .B2(n3403), .C1(n2530), 
        .C2(n6834), .ZN(n6048) );
  inv0d0 U3490 ( .I(debug_bus_rsp_data[25]), .ZN(n2512) );
  aoi22d1 U3491 ( .A1(iBus_rsp_payload_data[25]), .A2(n2523), .B1(
        writeBack_REGFILE_WRITE_DATA[25]), .B2(n2522), .ZN(n2511) );
  nd02d0 U3492 ( .A1(n2529), .A2(n2511), .ZN(n3259) );
  inv0d0 U3493 ( .I(n3259), .ZN(n3402) );
  inv0d0 U3494 ( .I(execute_PC[25]), .ZN(n6829) );
  oai222d1 U3495 ( .A1(n2512), .A2(n2514), .B1(n2531), .B2(n3402), .C1(n2530), 
        .C2(n6829), .ZN(n6047) );
  inv0d0 U3496 ( .I(debug_bus_rsp_data[26]), .ZN(n2515) );
  aoi22d1 U3497 ( .A1(iBus_rsp_payload_data[26]), .A2(n2523), .B1(
        writeBack_REGFILE_WRITE_DATA[26]), .B2(n2522), .ZN(n2513) );
  nd02d0 U3498 ( .A1(n2529), .A2(n2513), .ZN(n3258) );
  inv0d0 U3499 ( .I(n3258), .ZN(n3401) );
  inv0d0 U3500 ( .I(execute_PC[26]), .ZN(n6824) );
  oai222d1 U3501 ( .A1(n2515), .A2(n2514), .B1(n2531), .B2(n3401), .C1(n2530), 
        .C2(n6824), .ZN(n6046) );
  inv0d0 U3502 ( .I(debug_bus_rsp_data[27]), .ZN(n2517) );
  aoi22d1 U3503 ( .A1(iBus_rsp_payload_data[27]), .A2(n2523), .B1(
        writeBack_REGFILE_WRITE_DATA[27]), .B2(n2522), .ZN(n2516) );
  nd02d0 U3504 ( .A1(n2529), .A2(n2516), .ZN(n3257) );
  inv0d0 U3505 ( .I(n3257), .ZN(n3400) );
  inv0d0 U3506 ( .I(execute_PC[27]), .ZN(n6819) );
  oai222d1 U3507 ( .A1(n2517), .A2(n2532), .B1(n2531), .B2(n3400), .C1(n2530), 
        .C2(n6819), .ZN(n6045) );
  inv0d0 U3508 ( .I(debug_bus_rsp_data[28]), .ZN(n2519) );
  aoi22d1 U3509 ( .A1(iBus_rsp_payload_data[28]), .A2(n2523), .B1(
        writeBack_REGFILE_WRITE_DATA[28]), .B2(n2522), .ZN(n2518) );
  nd02d0 U3510 ( .A1(n2529), .A2(n2518), .ZN(n3256) );
  inv0d0 U3511 ( .I(n3256), .ZN(n3399) );
  inv0d0 U3512 ( .I(execute_PC[28]), .ZN(n6814) );
  oai222d1 U3513 ( .A1(n2519), .A2(n2532), .B1(n2531), .B2(n3399), .C1(n2530), 
        .C2(n6814), .ZN(n6044) );
  inv0d0 U3514 ( .I(debug_bus_rsp_data[29]), .ZN(n2521) );
  aoi22d1 U3515 ( .A1(iBus_rsp_payload_data[29]), .A2(n2523), .B1(
        writeBack_REGFILE_WRITE_DATA[29]), .B2(n2522), .ZN(n2520) );
  nd02d0 U3516 ( .A1(n2529), .A2(n2520), .ZN(n3254) );
  inv0d0 U3517 ( .I(n3254), .ZN(n3397) );
  inv0d0 U3518 ( .I(execute_PC[29]), .ZN(n6809) );
  oai222d1 U3519 ( .A1(n2521), .A2(n2532), .B1(n2531), .B2(n3397), .C1(n2530), 
        .C2(n6809), .ZN(n6043) );
  inv0d0 U3520 ( .I(debug_bus_rsp_data[30]), .ZN(n2525) );
  aoi22d1 U3521 ( .A1(iBus_rsp_payload_data[30]), .A2(n2523), .B1(
        writeBack_REGFILE_WRITE_DATA[30]), .B2(n2522), .ZN(n2524) );
  nd02d0 U3522 ( .A1(n2529), .A2(n2524), .ZN(n3253) );
  inv0d0 U3523 ( .I(n3253), .ZN(n3396) );
  inv0d0 U3524 ( .I(execute_PC[30]), .ZN(n6418) );
  oai222d1 U3525 ( .A1(n2525), .A2(n2532), .B1(n2531), .B2(n3396), .C1(n2530), 
        .C2(n6418), .ZN(n6042) );
  inv0d0 U3526 ( .I(debug_bus_rsp_data[31]), .ZN(n2533) );
  aoi22d1 U3527 ( .A1(n2527), .A2(iBus_rsp_payload_data[31]), .B1(
        writeBack_REGFILE_WRITE_DATA[31]), .B2(n2526), .ZN(n2528) );
  nd02d0 U3528 ( .A1(n2529), .A2(n2528), .ZN(n3252) );
  inv0d0 U3529 ( .I(n3252), .ZN(n3395) );
  inv0d0 U3530 ( .I(execute_PC[31]), .ZN(n6416) );
  oai222d1 U3531 ( .A1(n2533), .A2(n2532), .B1(n2531), .B2(n3395), .C1(n2530), 
        .C2(n6416), .ZN(n6041) );
  oaim21d1 U3532 ( .B1(n3673), .B2(CsrPlugin_mcause_interrupt), .A(n2534), 
        .ZN(n6040) );
  mx02d1 U3533 ( .I0(CsrPlugin_mtval[0]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[0]), .S(n3671), 
        .Z(n6039) );
  mx02d1 U3534 ( .I0(CsrPlugin_mtval[31]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[31]), .S(n3671), 
        .Z(n6038) );
  mx02d1 U3535 ( .I0(CsrPlugin_mtval[30]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[30]), .S(n3671), 
        .Z(n6037) );
  mx02d1 U3536 ( .I0(CsrPlugin_mtval[29]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[29]), .S(n3671), 
        .Z(n6036) );
  inv0d1 U3537 ( .I(n3673), .ZN(n3676) );
  mx02d1 U3538 ( .I0(CsrPlugin_mtval[28]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[28]), .S(n3676), 
        .Z(n6035) );
  mx02d1 U3539 ( .I0(CsrPlugin_mtval[27]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[27]), .S(n3676), 
        .Z(n6034) );
  mx02d1 U3540 ( .I0(CsrPlugin_mtval[26]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[26]), .S(n3676), 
        .Z(n6033) );
  mx02d1 U3541 ( .I0(CsrPlugin_mtval[25]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[25]), .S(n3676), 
        .Z(n6032) );
  mx02d1 U3542 ( .I0(CsrPlugin_mtval[24]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[24]), .S(n3676), 
        .Z(n6031) );
  mx02d1 U3543 ( .I0(CsrPlugin_mtval[23]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[23]), .S(n3676), 
        .Z(n6030) );
  mx02d1 U3544 ( .I0(CsrPlugin_mtval[22]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[22]), .S(n3676), 
        .Z(n6029) );
  mx02d1 U3545 ( .I0(CsrPlugin_mtval[21]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[21]), .S(n3676), 
        .Z(n6028) );
  mx02d1 U3546 ( .I0(CsrPlugin_mtval[20]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[20]), .S(n3676), 
        .Z(n6027) );
  mx02d1 U3547 ( .I0(CsrPlugin_mtval[19]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[19]), .S(
        CsrPlugin_hadException), .Z(n6026) );
  mx02d1 U3548 ( .I0(CsrPlugin_mtval[18]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[18]), .S(
        CsrPlugin_hadException), .Z(n6025) );
  mx02d1 U3549 ( .I0(CsrPlugin_mtval[17]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[17]), .S(
        CsrPlugin_hadException), .Z(n6024) );
  mx02d1 U3550 ( .I0(CsrPlugin_mtval[16]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[16]), .S(
        CsrPlugin_hadException), .Z(n6023) );
  mx02d1 U3551 ( .I0(CsrPlugin_mtval[15]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[15]), .S(
        CsrPlugin_hadException), .Z(n6022) );
  mx02d1 U3552 ( .I0(CsrPlugin_mtval[14]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[14]), .S(
        CsrPlugin_hadException), .Z(n6021) );
  mx02d1 U3553 ( .I0(CsrPlugin_mtval[13]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[13]), .S(
        CsrPlugin_hadException), .Z(n6020) );
  mx02d1 U3554 ( .I0(CsrPlugin_mtval[12]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[12]), .S(
        CsrPlugin_hadException), .Z(n6019) );
  mx02d1 U3555 ( .I0(CsrPlugin_mtval[11]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[11]), .S(n3676), 
        .Z(n6018) );
  mx02d1 U3556 ( .I0(CsrPlugin_mtval[10]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[10]), .S(
        CsrPlugin_hadException), .Z(n6017) );
  mx02d1 U3557 ( .I0(CsrPlugin_mtval[9]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[9]), .S(n3676), 
        .Z(n6016) );
  mx02d1 U3558 ( .I0(CsrPlugin_mtval[8]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[8]), .S(
        CsrPlugin_hadException), .Z(n6015) );
  mx02d1 U3559 ( .I0(CsrPlugin_mtval[7]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[7]), .S(
        CsrPlugin_hadException), .Z(n6014) );
  mx02d1 U3560 ( .I0(CsrPlugin_mtval[6]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[6]), .S(n3676), 
        .Z(n6013) );
  mx02d1 U3561 ( .I0(CsrPlugin_mtval[5]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[5]), .S(
        CsrPlugin_hadException), .Z(n6012) );
  mx02d1 U3562 ( .I0(CsrPlugin_mtval[4]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[4]), .S(n3676), 
        .Z(n6011) );
  mx02d1 U3563 ( .I0(CsrPlugin_mtval[3]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[3]), .S(
        CsrPlugin_hadException), .Z(n6010) );
  aoim22d1 U3564 ( .A1(n2535), .A2(n3673), .B1(n3673), .B2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[2]), .Z(n6009) );
  mx02d1 U3565 ( .I0(CsrPlugin_mtval[1]), .I1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr[1]), .S(n3676), 
        .Z(n6008) );
  mx02d1 U3566 ( .I0(execute_RS2[0]), .I1(_zz_RegFilePlugin_regFile_port1[0]), 
        .S(n3558), .Z(n6007) );
  inv0d1 U3567 ( .I(n3232), .ZN(n3209) );
  oai22d1 U3568 ( .A1(n3209), .A2(n2537), .B1(n2536), .B2(n2605), .ZN(n6006)
         );
  nd04d0 U3569 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13[28]), .A2(
        _zz_decode_LEGAL_INSTRUCTION_13[29]), .A3(n2543), .A4(n2615), .ZN(
        n2549) );
  nd02d0 U3570 ( .A1(\_zz__zz_decode_ENV_CTRL_2_1[20] ), .A2(n2540), .ZN(n2542) );
  oai22d1 U3571 ( .A1(n2589), .A2(n2538), .B1(n2542), .B2(n2616), .ZN(n6005)
         );
  nr02d0 U3572 ( .A1(n2616), .A2(\_zz__zz_decode_ENV_CTRL_2_1[20] ), .ZN(n2539) );
  aor22d1 U3573 ( .A1(n3243), .A2(execute_CsrPlugin_csr_834), .B1(n2540), .B2(
        n2539), .Z(n6004) );
  oai22d1 U3574 ( .A1(decode_INSTRUCTION_21), .A2(n2542), .B1(n2589), .B2(
        n2541), .ZN(n6003) );
  inv0d0 U3575 ( .I(execute_CsrPlugin_csr_773), .ZN(n3560) );
  nd03d0 U3576 ( .A1(_zz_decode_LEGAL_INSTRUCTION_13[28]), .A2(
        _zz_decode_LEGAL_INSTRUCTION_13[29]), .A3(n2543), .ZN(n2544) );
  nr03d0 U3577 ( .A1(n3238), .A2(n2615), .A3(n2544), .ZN(n2547) );
  oai22d1 U3578 ( .A1(n2620), .A2(n3560), .B1(n2546), .B2(n2617), .ZN(n6002)
         );
  oai22d1 U3579 ( .A1(\_zz__zz_decode_ENV_CTRL_2_1[20] ), .A2(n2546), .B1(
        n2589), .B2(n2545), .ZN(n6001) );
  aor22d1 U3580 ( .A1(n2548), .A2(n2547), .B1(execute_CsrPlugin_csr_836), .B2(
        n3243), .Z(n6000) );
  oaim22d1 U3581 ( .A1(n2550), .A2(n2549), .B1(n3235), .B2(
        execute_CsrPlugin_csr_768), .ZN(n5999) );
  nd02d0 U3582 ( .A1(n3558), .A2(_zz_decode_LEGAL_INSTRUCTION_1_13), .ZN(n2626) );
  inv0d0 U3583 ( .I(n2626), .ZN(n2573) );
  aoi22d1 U3584 ( .A1(n2573), .A2(n2552), .B1(n3238), .B2(n2551), .ZN(n5998)
         );
  nr02d0 U3585 ( .A1(n3238), .A2(n2553), .ZN(n3045) );
  nr02d0 U3586 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1_13), .A2(n2554), .ZN(n2591) );
  inv0d0 U3587 ( .I(n2571), .ZN(n2568) );
  aoi31d1 U3588 ( .B1(_zz_decode_LEGAL_INSTRUCTION_1[5]), .B2(n3558), .B3(
        n2595), .A(n2568), .ZN(n2558) );
  inv0d0 U3589 ( .I(n2556), .ZN(n2582) );
  nd04d0 U3590 ( .A1(n2582), .A2(_zz_decode_LEGAL_INSTRUCTION_1[4]), .A3(
        decode_INSTRUCTION_30), .A4(n2625), .ZN(n2557) );
  aon211d1 U3591 ( .C1(n2577), .C2(n2586), .B(
        _zz_decode_LEGAL_INSTRUCTION_1[2]), .A(n2557), .ZN(n2593) );
  oai22d1 U3592 ( .A1(n2620), .A2(n2897), .B1(n2558), .B2(n2593), .ZN(n5997)
         );
  inv0d0 U3593 ( .I(execute_ENV_CTRL[0]), .ZN(n6801) );
  nd02d0 U3594 ( .A1(n3558), .A2(n2559), .ZN(n2561) );
  oai22d1 U3595 ( .A1(n2620), .A2(n6801), .B1(n2561), .B2(n2560), .ZN(n5996)
         );
  oaim22d1 U3596 ( .A1(n3209), .A2(n6802), .B1(n2617), .B2(n2562), .ZN(n5995)
         );
  aoim22d1 U3597 ( .A1(n3558), .A2(n2563), .B1(execute_IS_CSR), .B2(n3558), 
        .Z(n5994) );
  inv0d0 U3598 ( .I(execute_BRANCH_CTRL[0]), .ZN(n6268) );
  nd02d0 U3599 ( .A1(n2620), .A2(_zz_decode_LEGAL_INSTRUCTION_1[6]), .ZN(n2629) );
  inv0d0 U3600 ( .I(n2565), .ZN(n2564) );
  oai22d1 U3601 ( .A1(n3209), .A2(n6268), .B1(n2629), .B2(n2564), .ZN(n5993)
         );
  inv0d1 U3602 ( .I(n3247), .ZN(n3548) );
  inv0d0 U3603 ( .I(execute_BRANCH_CTRL[1]), .ZN(n6302) );
  nd03d0 U3604 ( .A1(n2589), .A2(_zz_decode_LEGAL_INSTRUCTION_1[2]), .A3(n2565), .ZN(n2567) );
  nd03d0 U3605 ( .A1(n2589), .A2(_zz_decode_LEGAL_INSTRUCTION_1[6]), .A3(
        _zz_decode_LEGAL_INSTRUCTION_1[3]), .ZN(n2566) );
  oai211d1 U3606 ( .C1(n3548), .C2(n6302), .A(n2567), .B(n2566), .ZN(n5992) );
  oai21d1 U3607 ( .B1(decode_INSTRUCTION_30), .B2(n2625), .A(n2568), .ZN(n2569) );
  oai21d1 U3608 ( .B1(n2589), .B2(n2570), .A(n2569), .ZN(n5991) );
  oai22d1 U3609 ( .A1(n2620), .A2(n2572), .B1(n2625), .B2(n2571), .ZN(n5990)
         );
  nd02d0 U3610 ( .A1(n3209), .A2(_zz_decode_LEGAL_INSTRUCTION_7_12), .ZN(n2574) );
  aor22d1 U3611 ( .A1(n2621), .A2(execute_ALU_BITWISE_CTRL[0]), .B1(n2574), 
        .B2(n2573), .Z(n5989) );
  oai21d1 U3612 ( .B1(n3558), .B2(n6681), .A(n2574), .ZN(n5988) );
  inv0d0 U3613 ( .I(execute_SRC_LESS_UNSIGNED), .ZN(n2636) );
  oai222d1 U3614 ( .A1(n2636), .A2(n3558), .B1(n2626), .B2(
        _zz_decode_LEGAL_INSTRUCTION_1[4]), .C1(n2574), .C2(
        \_zz_decode_LEGAL_INSTRUCTION_7[14] ), .ZN(n5987) );
  aoi221d1 U3615 ( .B1(_zz_decode_LEGAL_INSTRUCTION_1[3]), .B2(n2577), .C1(
        n2575), .C2(n2582), .A(n3238), .ZN(n2576) );
  oan211d1 U3616 ( .C1(n2578), .C2(n2577), .B(n3045), .A(n2576), .ZN(n2579) );
  inv0d0 U3617 ( .I(execute_REGFILE_WRITE_VALID), .ZN(n6804) );
  oai22d1 U3618 ( .A1(n2580), .A2(n2579), .B1(n2589), .B2(n6804), .ZN(n5986)
         );
  aoi22d1 U3619 ( .A1(n3209), .A2(n2582), .B1(n2581), .B2(n2621), .ZN(n5985)
         );
  nr02d0 U3620 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[6]), .A2(
        _zz_decode_LEGAL_INSTRUCTION_1[4]), .ZN(n2592) );
  inv0d1 U3621 ( .I(n3238), .ZN(n3516) );
  aon211d1 U3622 ( .C1(_zz_decode_LEGAL_INSTRUCTION_1[5]), .C2(n2592), .B(
        _zz_decode_LEGAL_INSTRUCTION_1[2]), .A(n3516), .ZN(n2583) );
  oai21d1 U3623 ( .B1(n2589), .B2(n2584), .A(n2583), .ZN(n5984) );
  inv0d1 U3624 ( .I(n3232), .ZN(n3249) );
  nd02d0 U3625 ( .A1(n3249), .A2(n2585), .ZN(n2587) );
  oai22d1 U3626 ( .A1(n2620), .A2(n2588), .B1(n2587), .B2(n2586), .ZN(n5983)
         );
  nd03d0 U3627 ( .A1(\_zz_decode_LEGAL_INSTRUCTION_7[14] ), .A2(n3045), .A3(
        n3047), .ZN(n2590) );
  inv0d0 U3628 ( .I(execute_ALU_CTRL[1]), .ZN(n2639) );
  oai22d1 U3629 ( .A1(n2591), .A2(n2590), .B1(n2589), .B2(n2639), .ZN(n5982)
         );
  nr02d0 U3630 ( .A1(n3238), .A2(_zz_decode_LEGAL_INSTRUCTION_1[3]), .ZN(n3046) );
  aor22d1 U3631 ( .A1(n3243), .A2(execute_MEMORY_ENABLE), .B1(n3046), .B2(
        n2592), .Z(n5981) );
  aoim22d1 U3632 ( .A1(n2594), .A2(n3243), .B1(n3238), .B2(n2593), .Z(n5980)
         );
  nd02d0 U3633 ( .A1(n3558), .A2(n2595), .ZN(n2596) );
  nd03d0 U3634 ( .A1(_zz_decode_LEGAL_INSTRUCTION_1[6]), .A2(
        \_zz_decode_LEGAL_INSTRUCTION_7[14] ), .A3(n3045), .ZN(n2599) );
  oai211d1 U3635 ( .C1(n3516), .C2(n2597), .A(n2596), .B(n2599), .ZN(n5979) );
  inv0d1 U3636 ( .I(n3238), .ZN(n3526) );
  inv0d1 U3637 ( .I(n3232), .ZN(n3559) );
  nd02d0 U3638 ( .A1(n3559), .A2(n2598), .ZN(n2600) );
  oai211d1 U3639 ( .C1(n3526), .C2(n2601), .A(n2600), .B(n2599), .ZN(n5978) );
  oai22d1 U3640 ( .A1(n2621), .A2(_zz_decode_LEGAL_INSTRUCTION_1[0]), .B1(
        execute_INSTRUCTION[0]), .B2(n3558), .ZN(n2602) );
  inv0d0 U3641 ( .I(n2602), .ZN(n5977) );
  aoi22d1 U3642 ( .A1(n2620), .A2(n2603), .B1(n6284), .B2(n2621), .ZN(n5976)
         );
  aoi22d1 U3643 ( .A1(n2620), .A2(n2605), .B1(n2604), .B2(n2621), .ZN(n5975)
         );
  aoim22d1 U3644 ( .A1(n6459), .A2(n3243), .B1(n3243), .B2(
        _zz_decode_LEGAL_INSTRUCTION_13[29]), .Z(n5974) );
  aoi22d1 U3645 ( .A1(n2620), .A2(n2606), .B1(n6474), .B2(n2621), .ZN(n5973)
         );
  aoi22d1 U3646 ( .A1(n2620), .A2(n2608), .B1(n2607), .B2(n2621), .ZN(n5972)
         );
  aoi22d1 U3647 ( .A1(n2620), .A2(n2610), .B1(n2609), .B2(n2621), .ZN(n5971)
         );
  aoi22d1 U3648 ( .A1(n2620), .A2(n2612), .B1(n2611), .B2(n2621), .ZN(n5970)
         );
  aoi22d1 U3649 ( .A1(n2620), .A2(n2613), .B1(n6293), .B2(n2621), .ZN(n5969)
         );
  aoi22d1 U3650 ( .A1(n2620), .A2(n2614), .B1(n6295), .B2(n3247), .ZN(n5968)
         );
  aoi22d1 U3651 ( .A1(n3209), .A2(n2615), .B1(n6298), .B2(n2621), .ZN(n5967)
         );
  aoi22d1 U3652 ( .A1(n2620), .A2(n2616), .B1(n6303), .B2(n2621), .ZN(n5966)
         );
  aoi22d1 U3653 ( .A1(n2620), .A2(n2617), .B1(n6307), .B2(n3247), .ZN(n5965)
         );
  aoi22d1 U3654 ( .A1(n3209), .A2(n2618), .B1(n6269), .B2(n2621), .ZN(n5964)
         );
  aoi22d1 U3655 ( .A1(n2620), .A2(n173), .B1(n6271), .B2(n2621), .ZN(n5963) );
  inv0d0 U3656 ( .I(_zz__zz_execute_SRC1_1[2]), .ZN(n6273) );
  aoi22d1 U3657 ( .A1(n3209), .A2(n2622), .B1(n6273), .B2(n2621), .ZN(n5962)
         );
  aoi22d1 U3658 ( .A1(n3209), .A2(n2623), .B1(n6275), .B2(n3247), .ZN(n5961)
         );
  aoi22d1 U3659 ( .A1(n3209), .A2(n174), .B1(n6277), .B2(n3247), .ZN(n5960) );
  aoi22d1 U3660 ( .A1(n3209), .A2(n2625), .B1(n6650), .B2(n3247), .ZN(n5959)
         );
  oai21d1 U3661 ( .B1(n3558), .B2(n6919), .A(n2626), .ZN(n5958) );
  inv0d0 U3662 ( .I(_zz__zz_execute_SRC2_3[4]), .ZN(n6694) );
  aoi22d1 U3663 ( .A1(n3209), .A2(n2627), .B1(n6694), .B2(n3247), .ZN(n5957)
         );
  aoi22d1 U3664 ( .A1(n3209), .A2(n2628), .B1(n6709), .B2(n3247), .ZN(n5956)
         );
  aoim22d1 U3665 ( .A1(n6722), .A2(n3238), .B1(n3238), .B2(
        decode_INSTRUCTION_9), .Z(n5955) );
  aoim22d1 U3666 ( .A1(n6753), .A2(n3243), .B1(n3238), .B2(
        decode_INSTRUCTION_7), .Z(n5953) );
  oaim21d1 U3667 ( .B1(n3235), .B2(execute_INSTRUCTION[6]), .A(n2629), .ZN(
        n5952) );
  aoi22d1 U3668 ( .A1(n3209), .A2(n2630), .B1(n6781), .B2(n3232), .ZN(n5951)
         );
  aoi22d1 U3669 ( .A1(memory_REGFILE_WRITE_DATA[1]), .A2(n3027), .B1(n2870), 
        .B2(n3039), .ZN(n2648) );
  nr02d0 U3670 ( .A1(n3036), .A2(n2631), .ZN(n2632) );
  aoi22d1 U3671 ( .A1(n3036), .A2(n2631), .B1(n3678), .B2(n2644), .ZN(n3752)
         );
  aoi22d1 U3672 ( .A1(n2761), .A2(n2632), .B1(n2960), .B2(n3752), .ZN(n2642)
         );
  inv0d0 U3673 ( .I(n6805), .ZN(n2634) );
  oai22d1 U3674 ( .A1(n2634), .A2(n3754), .B1(n2636), .B2(n2633), .ZN(n2635)
         );
  aoi31d1 U3675 ( .B1(n2638), .B2(n2637), .B3(n2636), .A(n2635), .ZN(n3782) );
  nd04d0 U3676 ( .A1(execute_ALU_CTRL[0]), .A2(n3782), .A3(n2640), .A4(n2639), 
        .ZN(n2641) );
  oai211d1 U3677 ( .C1(n3025), .C2(n6994), .A(n2642), .B(n2641), .ZN(n2643) );
  oan211d1 U3678 ( .C1(n3678), .C2(n2644), .B(n3026), .A(n2643), .ZN(n2647) );
  aoi22d1 U3679 ( .A1(n2872), .A2(n2645), .B1(memory_REGFILE_WRITE_DATA[0]), 
        .B2(n299), .ZN(n2646) );
  aon211d1 U3680 ( .C1(n2648), .C2(n2647), .B(n2996), .A(n2646), .ZN(n5950) );
  aoi22d1 U3681 ( .A1(memory_REGFILE_WRITE_DATA[29]), .A2(n2984), .B1(n2870), 
        .B2(n2649), .ZN(n2663) );
  aoi22d1 U3682 ( .A1(execute_SRC2_FORCE_ZERO), .A2(n2659), .B1(n2652), .B2(
        n2897), .ZN(n6806) );
  aoi22d1 U3683 ( .A1(n2761), .A2(n2654), .B1(n2969), .B2(n2670), .ZN(n2656)
         );
  mx02d1 U3684 ( .I0(n2659), .I1(n2671), .S(n2658), .Z(n3743) );
  aoi22d1 U3685 ( .A1(n2818), .A2(memory_REGFILE_WRITE_DATA[31]), .B1(n2960), 
        .B2(n3743), .ZN(n2655) );
  oai211d1 U3686 ( .C1(n3025), .C2(n6806), .A(n2656), .B(n2655), .ZN(n2657) );
  oan211d1 U3687 ( .C1(n2659), .C2(n2658), .B(n3026), .A(n2657), .ZN(n2662) );
  aoi22d1 U3688 ( .A1(n2872), .A2(n2660), .B1(memory_REGFILE_WRITE_DATA[30]), 
        .B2(n299), .ZN(n2661) );
  aon211d1 U3689 ( .C1(n2663), .C2(n2662), .B(n2996), .A(n2661), .ZN(n5949) );
  aoi22d1 U3690 ( .A1(n2872), .A2(n2664), .B1(n2989), .B2(n2665), .ZN(n2678)
         );
  aoi22d1 U3691 ( .A1(n3026), .A2(n2670), .B1(n2969), .B2(n2694), .ZN(n2676)
         );
  aoi22d1 U3692 ( .A1(n3027), .A2(memory_REGFILE_WRITE_DATA[30]), .B1(n3029), 
        .B2(memory_REGFILE_WRITE_DATA[28]), .ZN(n2675) );
  mx02d1 U3693 ( .I0(n2670), .I1(n2682), .S(n2665), .Z(n3762) );
  aoi22d1 U3694 ( .A1(execute_SRC2_FORCE_ZERO), .A2(n2670), .B1(n2669), .B2(
        n2897), .ZN(n6811) );
  oai22d1 U3695 ( .A1(n2671), .A2(n314), .B1(n3025), .B2(n6811), .ZN(n2672) );
  aoi211d1 U3696 ( .C1(n3762), .C2(n3032), .A(n2673), .B(n2672), .ZN(n2674) );
  aor31d1 U3697 ( .B1(n2676), .B2(n2675), .B3(n2674), .A(n2996), .Z(n2677) );
  oaim211d1 U3698 ( .C1(n299), .C2(memory_REGFILE_WRITE_DATA[29]), .A(n2678), 
        .B(n2677), .ZN(n5948) );
  aoi22d1 U3699 ( .A1(execute_SRC2_FORCE_ZERO), .A2(n2694), .B1(n2681), .B2(
        n2897), .ZN(n6816) );
  oai22d1 U3700 ( .A1(n2682), .A2(n314), .B1(n3025), .B2(n6816), .ZN(n2687) );
  mx02d1 U3701 ( .I0(n2694), .I1(n2683), .S(n2689), .Z(n3758) );
  aoi22d1 U3702 ( .A1(n2818), .A2(memory_REGFILE_WRITE_DATA[29]), .B1(n2960), 
        .B2(n3758), .ZN(n2685) );
  aon211d1 U3703 ( .C1(n2761), .C2(n2689), .B(n3026), .A(n2694), .ZN(n2684) );
  nd02d0 U3704 ( .A1(n2685), .A2(n2684), .ZN(n2686) );
  aoi211d1 U3705 ( .C1(n2984), .C2(memory_REGFILE_WRITE_DATA[27]), .A(n2687), 
        .B(n2686), .ZN(n2692) );
  aoi22d1 U3706 ( .A1(n2872), .A2(n2688), .B1(memory_REGFILE_WRITE_DATA[28]), 
        .B2(n299), .ZN(n2691) );
  aoi22d1 U3707 ( .A1(n2989), .A2(n2689), .B1(n2923), .B2(n2711), .ZN(n2690)
         );
  oai211d1 U3708 ( .C1(n2692), .C2(n2996), .A(n2691), .B(n2690), .ZN(n5947) );
  aoi22d1 U3709 ( .A1(n2999), .A2(n2693), .B1(n2989), .B2(n2695), .ZN(n2707)
         );
  aoi22d1 U3710 ( .A1(n3026), .A2(n2711), .B1(n3029), .B2(
        memory_REGFILE_WRITE_DATA[26]), .ZN(n2705) );
  aoi22d1 U3711 ( .A1(n2870), .A2(n2694), .B1(n2969), .B2(n2713), .ZN(n2704)
         );
  mx02d1 U3712 ( .I0(n2711), .I1(n2697), .S(n2695), .Z(n3742) );
  nr03d0 U3713 ( .A1(n2697), .A2(n2696), .A3(n2961), .ZN(n2702) );
  aoi22d1 U3714 ( .A1(execute_SRC2_FORCE_ZERO), .A2(n2711), .B1(n2700), .B2(
        n2897), .ZN(n6821) );
  oaim22d1 U3715 ( .A1(n3005), .A2(n6821), .B1(n2818), .B2(
        memory_REGFILE_WRITE_DATA[28]), .ZN(n2701) );
  aoi211d1 U3716 ( .C1(n3742), .C2(n3032), .A(n2702), .B(n2701), .ZN(n2703) );
  aor31d1 U3717 ( .B1(n2705), .B2(n2704), .B3(n2703), .A(n3033), .Z(n2706) );
  oaim211d1 U3718 ( .C1(n299), .C2(memory_REGFILE_WRITE_DATA[27]), .A(n2707), 
        .B(n2706), .ZN(n5946) );
  aoi22d1 U3719 ( .A1(execute_SRC2_FORCE_ZERO), .A2(n2713), .B1(n2710), .B2(
        n2897), .ZN(n6826) );
  mx02d1 U3720 ( .I0(n2713), .I1(n2724), .S(n2712), .Z(n3737) );
  oaim22d1 U3721 ( .A1(n3005), .A2(n6826), .B1(n3032), .B2(n3737), .ZN(n2718)
         );
  aoi22d1 U3722 ( .A1(n3026), .A2(n2713), .B1(n2870), .B2(n2711), .ZN(n2716)
         );
  aoi22d1 U3723 ( .A1(n2969), .A2(n2728), .B1(n3029), .B2(
        memory_REGFILE_WRITE_DATA[25]), .ZN(n2715) );
  aon211d1 U3724 ( .C1(n2761), .C2(n2713), .B(n3026), .A(n2712), .ZN(n2714) );
  aoi211d1 U3725 ( .C1(n3027), .C2(memory_REGFILE_WRITE_DATA[27]), .A(n2718), 
        .B(n2717), .ZN(n2720) );
  inv0d0 U3726 ( .I(memory_REGFILE_WRITE_DATA[26]), .ZN(n2723) );
  oai222d1 U3727 ( .A1(n3033), .A2(n2720), .B1(n2723), .B2(n2749), .C1(n2748), 
        .C2(n2719), .ZN(n5945) );
  nr02d0 U3728 ( .A1(n2739), .A2(n2721), .ZN(n3748) );
  oan211d1 U3729 ( .C1(n3748), .C2(n3013), .B(n3006), .A(n3749), .ZN(n2732) );
  oai22d1 U3730 ( .A1(n2724), .A2(n314), .B1(n2980), .B2(n2723), .ZN(n2731) );
  aoi22d1 U3731 ( .A1(execute_SRC2_FORCE_ZERO), .A2(n2728), .B1(n2727), .B2(
        n2897), .ZN(n6831) );
  oai22d1 U3732 ( .A1(n2754), .A2(n3035), .B1(n3025), .B2(n6831), .ZN(n2730)
         );
  inv0d0 U3733 ( .I(memory_REGFILE_WRITE_DATA[24]), .ZN(n2753) );
  oaim22d1 U3734 ( .A1(n2943), .A2(n2753), .B1(n2761), .B2(n3748), .ZN(n2729)
         );
  inv0d0 U3735 ( .I(memory_REGFILE_WRITE_DATA[25]), .ZN(n2734) );
  oai222d1 U3736 ( .A1(n3033), .A2(n2735), .B1(n2734), .B2(n2942), .C1(n2748), 
        .C2(n2733), .ZN(n5944) );
  aoi22d1 U3737 ( .A1(n2932), .A2(n2740), .B1(n2738), .B2(n2897), .ZN(n6836)
         );
  oai22d1 U3738 ( .A1(n2739), .A2(n314), .B1(n3005), .B2(n6836), .ZN(n2746) );
  aoi22d1 U3739 ( .A1(n2818), .A2(memory_REGFILE_WRITE_DATA[25]), .B1(n2969), 
        .B2(n2760), .ZN(n2744) );
  mx02d1 U3740 ( .I0(n2740), .I1(n2754), .S(n2741), .Z(n3736) );
  aoi22d1 U3741 ( .A1(n3026), .A2(n2741), .B1(n2960), .B2(n3736), .ZN(n2743)
         );
  aon211d1 U3742 ( .C1(n2761), .C2(n2741), .B(n3026), .A(n2740), .ZN(n2742) );
  aoi211d1 U3743 ( .C1(n3029), .C2(memory_REGFILE_WRITE_DATA[23]), .A(n2746), 
        .B(n2745), .ZN(n2750) );
  oai222d1 U3744 ( .A1(n3033), .A2(n2750), .B1(n2753), .B2(n2749), .C1(n2748), 
        .C2(n2747), .ZN(n5943) );
  aoi22d1 U3745 ( .A1(n2872), .A2(n2751), .B1(n2989), .B2(n2759), .ZN(n2769)
         );
  oai22d1 U3746 ( .A1(n2755), .A2(n3006), .B1(n2752), .B2(n3035), .ZN(n2767)
         );
  oai22d1 U3747 ( .A1(n2754), .A2(n314), .B1(n2980), .B2(n2753), .ZN(n2766) );
  mx02d1 U3748 ( .I0(n2760), .I1(n2755), .S(n2759), .Z(n3765) );
  aoi22d1 U3749 ( .A1(n2932), .A2(n2760), .B1(n2758), .B2(n2897), .ZN(n6841)
         );
  aoim22d1 U3750 ( .A1(n2960), .A2(n3765), .B1(n3005), .B2(n6841), .Z(n2763)
         );
  oai211d1 U3751 ( .C1(n2764), .C2(n2943), .A(n2763), .B(n2762), .ZN(n2765) );
  oai31d1 U3752 ( .B1(n2767), .B2(n2766), .B3(n2765), .A(n2856), .ZN(n2768) );
  oaim211d1 U3753 ( .C1(n299), .C2(memory_REGFILE_WRITE_DATA[23]), .A(n2769), 
        .B(n2768), .ZN(n5942) );
  inv0d0 U3754 ( .I(n2989), .ZN(n3043) );
  aoi22d1 U3755 ( .A1(n2872), .A2(n2770), .B1(memory_REGFILE_WRITE_DATA[21]), 
        .B2(n3020), .ZN(n2784) );
  mx02d1 U3756 ( .I0(n2782), .I1(n2790), .S(n2781), .Z(n3744) );
  aoi22d1 U3757 ( .A1(n2932), .A2(n2782), .B1(n2773), .B2(n2897), .ZN(n6851)
         );
  oai22d1 U3758 ( .A1(n2774), .A2(n3006), .B1(n3025), .B2(n6851), .ZN(n2778)
         );
  inv0d0 U3759 ( .I(memory_REGFILE_WRITE_DATA[20]), .ZN(n2804) );
  aoi22d1 U3760 ( .A1(n2870), .A2(n2775), .B1(n3027), .B2(
        memory_REGFILE_WRITE_DATA[22]), .ZN(n2776) );
  oai21d1 U3761 ( .B1(n2943), .B2(n2804), .A(n2776), .ZN(n2777) );
  aoi211d1 U3762 ( .C1(n3032), .C2(n3744), .A(n2778), .B(n2777), .ZN(n2779) );
  oan211d1 U3763 ( .C1(n2786), .C2(n3035), .B(n2779), .A(n2996), .ZN(n2780) );
  aoi31d1 U3764 ( .B1(n3040), .B2(n2782), .B3(n2781), .A(n2780), .ZN(n2783) );
  oai211d1 U3765 ( .C1(n2790), .C2(n3043), .A(n2784), .B(n2783), .ZN(n5940) );
  aoi22d1 U3766 ( .A1(n2999), .A2(n2785), .B1(n2989), .B2(n2805), .ZN(n2799)
         );
  mx02d1 U3767 ( .I0(n2805), .I1(n2786), .S(n2797), .Z(n3759) );
  aoi22d1 U3768 ( .A1(n2932), .A2(n2805), .B1(n2789), .B2(n2897), .ZN(n6856)
         );
  oai22d1 U3769 ( .A1(n2790), .A2(n314), .B1(n3025), .B2(n6856), .ZN(n2794) );
  aoi22d1 U3770 ( .A1(n3027), .A2(memory_REGFILE_WRITE_DATA[21]), .B1(n3029), 
        .B2(memory_REGFILE_WRITE_DATA[19]), .ZN(n2791) );
  oai21d1 U3771 ( .B1(n2792), .B2(n3006), .A(n2791), .ZN(n2793) );
  aoi211d1 U3772 ( .C1(n3032), .C2(n3759), .A(n2794), .B(n2793), .ZN(n2795) );
  oan211d1 U3773 ( .C1(n2819), .C2(n3035), .B(n2795), .A(n3033), .ZN(n2796) );
  aoi31d1 U3774 ( .B1(n3040), .B2(n2805), .B3(n2797), .A(n2796), .ZN(n2798) );
  oai211d1 U3775 ( .C1(n2942), .C2(n2804), .A(n2799), .B(n2798), .ZN(n5939) );
  aoi22d1 U3776 ( .A1(n2872), .A2(n2800), .B1(memory_REGFILE_WRITE_DATA[19]), 
        .B2(n3020), .ZN(n2814) );
  aoi22d1 U3777 ( .A1(n2932), .A2(n2812), .B1(n2803), .B2(n2897), .ZN(n6861)
         );
  oai22d1 U3778 ( .A1(n2980), .A2(n2804), .B1(n3025), .B2(n6861), .ZN(n2808)
         );
  inv0d0 U3779 ( .I(memory_REGFILE_WRITE_DATA[18]), .ZN(n2833) );
  mx02d1 U3780 ( .I0(n2812), .I1(n2819), .S(n2811), .Z(n3751) );
  aoi22d1 U3781 ( .A1(n2870), .A2(n2805), .B1(n2960), .B2(n3751), .ZN(n2806)
         );
  oai21d1 U3782 ( .B1(n2943), .B2(n2833), .A(n2806), .ZN(n2807) );
  aoi211d1 U3783 ( .C1(n3026), .C2(n2811), .A(n2808), .B(n2807), .ZN(n2809) );
  oan211d1 U3784 ( .C1(n2822), .C2(n3035), .B(n2809), .A(n2996), .ZN(n2810) );
  aoi31d1 U3785 ( .B1(n3040), .B2(n2812), .B3(n2811), .A(n2810), .ZN(n2813) );
  oai211d1 U3786 ( .C1(n2819), .C2(n3043), .A(n2814), .B(n2813), .ZN(n5938) );
  aoi22d1 U3787 ( .A1(n2932), .A2(n2835), .B1(n2817), .B2(n3003), .ZN(n6867)
         );
  oaim22d1 U3788 ( .A1(n3005), .A2(n6867), .B1(n2818), .B2(
        memory_REGFILE_WRITE_DATA[19]), .ZN(n2821) );
  oai22d1 U3789 ( .A1(n2822), .A2(n3006), .B1(n2819), .B2(n314), .ZN(n2820) );
  aoi211d1 U3790 ( .C1(n3029), .C2(memory_REGFILE_WRITE_DATA[17]), .A(n2821), 
        .B(n2820), .ZN(n2829) );
  mx02d1 U3791 ( .I0(n2835), .I1(n2822), .S(n2824), .Z(n3735) );
  aoi22d1 U3792 ( .A1(n2872), .A2(n2823), .B1(n2838), .B2(n2923), .ZN(n2826)
         );
  aon211d1 U3793 ( .C1(n3040), .C2(n2835), .B(n2989), .A(n2824), .ZN(n2825) );
  oai211d1 U3794 ( .C1(n2942), .C2(n2833), .A(n2826), .B(n2825), .ZN(n2827) );
  aoi21d1 U3795 ( .B1(n3735), .B2(n2994), .A(n2827), .ZN(n2828) );
  oai21d1 U3796 ( .B1(n2829), .B2(n2996), .A(n2828), .ZN(n5937) );
  aoi22d1 U3797 ( .A1(n2932), .A2(n2838), .B1(n2832), .B2(n3003), .ZN(n6872)
         );
  oai22d1 U3798 ( .A1(n6872), .A2(n3025), .B1(n2980), .B2(n2833), .ZN(n2834)
         );
  aoi21d1 U3799 ( .B1(n3029), .B2(memory_REGFILE_WRITE_DATA[16]), .A(n2834), 
        .ZN(n2846) );
  aoi22d1 U3800 ( .A1(n3026), .A2(n2839), .B1(n2870), .B2(n2835), .ZN(n2845)
         );
  mx02d1 U3801 ( .I0(n2838), .I1(n2836), .S(n2839), .Z(n3738) );
  inv0d0 U3802 ( .I(n2923), .ZN(n3019) );
  aoi22d1 U3803 ( .A1(n2872), .A2(n2837), .B1(memory_REGFILE_WRITE_DATA[17]), 
        .B2(n3020), .ZN(n2841) );
  aon211d1 U3804 ( .C1(n3040), .C2(n2839), .B(n2989), .A(n2838), .ZN(n2840) );
  oai211d1 U3805 ( .C1(n2842), .C2(n3019), .A(n2841), .B(n2840), .ZN(n2843) );
  aoi21d1 U3806 ( .B1(n2994), .B2(n3738), .A(n2843), .ZN(n2844) );
  aon211d1 U3807 ( .C1(n2846), .C2(n2845), .B(n2996), .A(n2844), .ZN(n5936) );
  aoi22d1 U3808 ( .A1(n2872), .A2(n2847), .B1(memory_REGFILE_WRITE_DATA[14]), 
        .B2(n3020), .ZN(n2859) );
  mx02d1 U3809 ( .I0(n2863), .I1(n2860), .S(n2862), .Z(n3773) );
  aoi22d1 U3810 ( .A1(n2870), .A2(n2848), .B1(n3029), .B2(
        memory_REGFILE_WRITE_DATA[13]), .ZN(n2854) );
  aoi22d1 U3811 ( .A1(n2932), .A2(n2863), .B1(n2851), .B2(n3003), .ZN(n6890)
         );
  oaim22d1 U3812 ( .A1(n3025), .A2(n6890), .B1(n3027), .B2(
        memory_REGFILE_WRITE_DATA[15]), .ZN(n2852) );
  aoi21d1 U3813 ( .B1(n3026), .B2(n2862), .A(n2852), .ZN(n2853) );
  oai211d1 U3814 ( .C1(n2855), .C2(n3035), .A(n2854), .B(n2853), .ZN(n2857) );
  aon211d1 U3815 ( .C1(n2960), .C2(n3773), .B(n2857), .A(n2856), .ZN(n2858) );
  oai211d1 U3816 ( .C1(n2860), .C2(n3043), .A(n2859), .B(n2858), .ZN(n2861) );
  aor31d1 U3817 ( .B1(n3040), .B2(n2863), .B3(n2862), .A(n2861), .Z(n5933) );
  aoi22d1 U3818 ( .A1(n2932), .A2(n2873), .B1(n2866), .B2(n3003), .ZN(n6902)
         );
  oai22d1 U3819 ( .A1(n6902), .A2(n3025), .B1(n2980), .B2(n2867), .ZN(n2868)
         );
  aoi21d1 U3820 ( .B1(n3026), .B2(n2874), .A(n2868), .ZN(n2880) );
  aoi22d1 U3821 ( .A1(n2870), .A2(n2869), .B1(n3029), .B2(
        memory_REGFILE_WRITE_DATA[10]), .ZN(n2879) );
  mx02d1 U3822 ( .I0(n2873), .I1(n2886), .S(n2874), .Z(n3739) );
  aoi22d1 U3823 ( .A1(n2872), .A2(n2871), .B1(memory_REGFILE_WRITE_DATA[11]), 
        .B2(n3020), .ZN(n2876) );
  aon211d1 U3824 ( .C1(n3040), .C2(n2874), .B(n2989), .A(n2873), .ZN(n2875) );
  oai211d1 U3825 ( .C1(n3019), .C2(n2900), .A(n2876), .B(n2875), .ZN(n2877) );
  aoi21d1 U3826 ( .B1(n2994), .B2(n3739), .A(n2877), .ZN(n2878) );
  aon211d1 U3827 ( .C1(n2880), .C2(n2879), .B(n3033), .A(n2878), .ZN(n5930) );
  aoi22d1 U3828 ( .A1(n2999), .A2(n2881), .B1(memory_REGFILE_WRITE_DATA[10]), 
        .B2(n3020), .ZN(n2894) );
  mx02d1 U3829 ( .I0(n2900), .I1(n2885), .S(n2890), .Z(n3761) );
  aoi22d1 U3830 ( .A1(n2932), .A2(n2885), .B1(n2884), .B2(n2897), .ZN(n6907)
         );
  oaim22d1 U3831 ( .A1(n6907), .A2(n3005), .B1(n3027), .B2(
        memory_REGFILE_WRITE_DATA[11]), .ZN(n2888) );
  inv0d0 U3832 ( .I(memory_REGFILE_WRITE_DATA[9]), .ZN(n2915) );
  oai22d1 U3833 ( .A1(n314), .A2(n2886), .B1(n2943), .B2(n2915), .ZN(n2887) );
  aoi211d1 U3834 ( .C1(n3032), .C2(n3761), .A(n2888), .B(n2887), .ZN(n2889) );
  oan211d1 U3835 ( .C1(n2890), .C2(n3006), .B(n2889), .A(n2996), .ZN(n2892) );
  inv0d0 U3836 ( .I(n3040), .ZN(n2927) );
  nr03d0 U3837 ( .A1(n2890), .A2(n2900), .A3(n2927), .ZN(n2891) );
  aoi211d1 U3838 ( .C1(n2923), .C2(n2899), .A(n2892), .B(n2891), .ZN(n2893) );
  oai211d1 U3839 ( .C1(n2900), .C2(n3043), .A(n2894), .B(n2893), .ZN(n5929) );
  mx02d1 U3840 ( .I0(n2916), .I1(n2899), .S(n2906), .Z(n3755) );
  aoi22d1 U3841 ( .A1(n2932), .A2(n2899), .B1(n2898), .B2(n2897), .ZN(n6913)
         );
  oaim22d1 U3842 ( .A1(n6913), .A2(n3005), .B1(n3027), .B2(
        memory_REGFILE_WRITE_DATA[10]), .ZN(n2902) );
  oai22d1 U3843 ( .A1(n2906), .A2(n3006), .B1(n314), .B2(n2900), .ZN(n2901) );
  aoi211d1 U3844 ( .C1(n3029), .C2(memory_REGFILE_WRITE_DATA[8]), .A(n2902), 
        .B(n2901), .ZN(n2903) );
  oan211d1 U3845 ( .C1(n3035), .C2(n2933), .B(n2903), .A(n2996), .ZN(n2908) );
  aoi22d1 U3846 ( .A1(n2999), .A2(n2904), .B1(memory_REGFILE_WRITE_DATA[9]), 
        .B2(n3020), .ZN(n2905) );
  oai31d1 U3847 ( .B1(n2906), .B2(n2916), .B3(n2927), .A(n2905), .ZN(n2907) );
  aoi211d1 U3848 ( .C1(n2994), .C2(n3755), .A(n2908), .B(n2907), .ZN(n2909) );
  oai21d1 U3849 ( .B1(n2916), .B2(n3043), .A(n2909), .ZN(n5928) );
  aoi22d1 U3850 ( .A1(n2999), .A2(n2910), .B1(memory_REGFILE_WRITE_DATA[8]), 
        .B2(n3020), .ZN(n2925) );
  mx02d1 U3851 ( .I0(n2933), .I1(n2914), .S(n2920), .Z(n3763) );
  aoi22d1 U3852 ( .A1(n2932), .A2(n2914), .B1(n2913), .B2(n3003), .ZN(n6918)
         );
  oai22d1 U3853 ( .A1(n6918), .A2(n3025), .B1(n2980), .B2(n2915), .ZN(n2918)
         );
  inv0d0 U3854 ( .I(memory_REGFILE_WRITE_DATA[7]), .ZN(n2944) );
  oai22d1 U3855 ( .A1(n314), .A2(n2916), .B1(n2943), .B2(n2944), .ZN(n2917) );
  aoi211d1 U3856 ( .C1(n3032), .C2(n3763), .A(n2918), .B(n2917), .ZN(n2919) );
  oan211d1 U3857 ( .C1(n2920), .C2(n3006), .B(n2919), .A(n2996), .ZN(n2922) );
  nr03d0 U3858 ( .A1(n2920), .A2(n2933), .A3(n2927), .ZN(n2921) );
  aoi211d1 U3859 ( .C1(n2923), .C2(n2931), .A(n2922), .B(n2921), .ZN(n2924) );
  oai211d1 U3860 ( .C1(n2933), .C2(n3043), .A(n2925), .B(n2924), .ZN(n5927) );
  aoi22d1 U3861 ( .A1(n2999), .A2(n2926), .B1(n2931), .B2(n2989), .ZN(n2941)
         );
  mx02d1 U3862 ( .I0(n2952), .I1(n2931), .S(n2934), .Z(n3750) );
  nr03d0 U3863 ( .A1(n2934), .A2(n2952), .A3(n2927), .ZN(n2939) );
  aoi22d1 U3864 ( .A1(n2932), .A2(n2931), .B1(n2930), .B2(n3003), .ZN(n6929)
         );
  oai22d1 U3865 ( .A1(n6929), .A2(n3025), .B1(n314), .B2(n2933), .ZN(n2936) );
  oaim22d1 U3866 ( .A1(n2934), .A2(n3006), .B1(n3027), .B2(
        memory_REGFILE_WRITE_DATA[8]), .ZN(n2935) );
  aoi211d1 U3867 ( .C1(n3029), .C2(memory_REGFILE_WRITE_DATA[6]), .A(n2936), 
        .B(n2935), .ZN(n2937) );
  oan211d1 U3868 ( .C1(n3035), .C2(n2966), .B(n2937), .A(n2996), .ZN(n2938) );
  aoi211d1 U3869 ( .C1(n2994), .C2(n3750), .A(n2939), .B(n2938), .ZN(n2940) );
  oai211d1 U3870 ( .C1(n2942), .C2(n2944), .A(n2941), .B(n2940), .ZN(n5926) );
  mx02d1 U3871 ( .I0(n2966), .I1(n2951), .S(n2947), .Z(n3760) );
  nr03d0 U3872 ( .A1(n2947), .A2(n2966), .A3(n2961), .ZN(n2946) );
  inv0d0 U3873 ( .I(memory_REGFILE_WRITE_DATA[5]), .ZN(n2979) );
  oai22d1 U3874 ( .A1(n2980), .A2(n2944), .B1(n2943), .B2(n2979), .ZN(n2945)
         );
  aoi211d1 U3875 ( .C1(n3760), .C2(n3032), .A(n2946), .B(n2945), .ZN(n2958) );
  aoi21d1 U3876 ( .B1(n2947), .B2(n2966), .A(n3006), .ZN(n2954) );
  aoi22d1 U3877 ( .A1(execute_SRC2_FORCE_ZERO), .A2(n2951), .B1(n2950), .B2(
        n3003), .ZN(n6943) );
  oai22d1 U3878 ( .A1(n6943), .A2(n3005), .B1(n314), .B2(n2952), .ZN(n2953) );
  aoi211d1 U3879 ( .C1(n2965), .C2(n2969), .A(n2954), .B(n2953), .ZN(n2957) );
  aoi22d1 U3880 ( .A1(n2999), .A2(n2955), .B1(memory_REGFILE_WRITE_DATA[6]), 
        .B2(n3020), .ZN(n2956) );
  aon211d1 U3881 ( .C1(n2958), .C2(n2957), .B(n2996), .A(n2956), .ZN(n5925) );
  aoi22d1 U3882 ( .A1(n2999), .A2(n2959), .B1(memory_REGFILE_WRITE_DATA[5]), 
        .B2(n3020), .ZN(n2974) );
  mx02d1 U3883 ( .I0(n2981), .I1(n2965), .S(n2975), .Z(n3764) );
  aoi22d1 U3884 ( .A1(n2984), .A2(memory_REGFILE_WRITE_DATA[4]), .B1(n2960), 
        .B2(n3764), .ZN(n2972) );
  aoi22d1 U3885 ( .A1(n3026), .A2(n2965), .B1(n3027), .B2(
        memory_REGFILE_WRITE_DATA[6]), .ZN(n2971) );
  aoi22d1 U3886 ( .A1(execute_SRC2_FORCE_ZERO), .A2(n2965), .B1(n2964), .B2(
        n3003), .ZN(n6949) );
  oai22d1 U3887 ( .A1(n6949), .A2(n3025), .B1(n314), .B2(n2966), .ZN(n2967) );
  aoi211d1 U3888 ( .C1(n2969), .C2(n2990), .A(n2968), .B(n2967), .ZN(n2970) );
  aor31d1 U3889 ( .B1(n2972), .B2(n2971), .B3(n2970), .A(n2996), .Z(n2973) );
  oai211d1 U3890 ( .C1(n2975), .C2(n3043), .A(n2974), .B(n2973), .ZN(n5924) );
  aoi22d1 U3891 ( .A1(execute_SRC2_FORCE_ZERO), .A2(n2990), .B1(n2978), .B2(
        n3003), .ZN(n6956) );
  oai22d1 U3892 ( .A1(n2980), .A2(n2979), .B1(n3005), .B2(n6956), .ZN(n2983)
         );
  oai22d1 U3893 ( .A1(n2985), .A2(n3006), .B1(n314), .B2(n2981), .ZN(n2982) );
  aoi211d1 U3894 ( .C1(n2984), .C2(memory_REGFILE_WRITE_DATA[3]), .A(n2983), 
        .B(n2982), .ZN(n2997) );
  aoi22d1 U3895 ( .A1(n2986), .A2(n2985), .B1(n2990), .B2(n2988), .ZN(n3734)
         );
  aoi22d1 U3896 ( .A1(n2999), .A2(n2987), .B1(memory_REGFILE_WRITE_DATA[4]), 
        .B2(n3020), .ZN(n2992) );
  aon211d1 U3897 ( .C1(n3040), .C2(n2990), .B(n2989), .A(n2988), .ZN(n2991) );
  oai211d1 U3898 ( .C1(n3008), .C2(n3019), .A(n2992), .B(n2991), .ZN(n2993) );
  aoi21d1 U3899 ( .B1(n3734), .B2(n2994), .A(n2993), .ZN(n2995) );
  oai21d1 U3900 ( .B1(n2997), .B2(n2996), .A(n2995), .ZN(n5923) );
  aoi22d1 U3901 ( .A1(n2999), .A2(n2998), .B1(memory_REGFILE_WRITE_DATA[2]), 
        .B2(n3020), .ZN(n3018) );
  aoi22d1 U3902 ( .A1(n3000), .A2(n3023), .B1(n3016), .B2(n3015), .ZN(n3772)
         );
  inv0d0 U3903 ( .I(n3772), .ZN(n3012) );
  aoi22d1 U3904 ( .A1(execute_SRC2_FORCE_ZERO), .A2(n3016), .B1(n3004), .B2(
        n3003), .ZN(n6973) );
  oaim22d1 U3905 ( .A1(n6973), .A2(n3005), .B1(n3027), .B2(
        memory_REGFILE_WRITE_DATA[3]), .ZN(n3010) );
  oai22d1 U3906 ( .A1(n3008), .A2(n314), .B1(n3007), .B2(n3006), .ZN(n3009) );
  aoi211d1 U3907 ( .C1(n3029), .C2(memory_REGFILE_WRITE_DATA[1]), .A(n3010), 
        .B(n3009), .ZN(n3011) );
  oan211d1 U3908 ( .C1(n3013), .C2(n3012), .B(n3011), .A(n3033), .ZN(n3014) );
  aoi31d1 U3909 ( .B1(n3016), .B2(n3040), .B3(n3015), .A(n3014), .ZN(n3017) );
  oai211d1 U3910 ( .C1(n3022), .C2(n3019), .A(n3018), .B(n3017), .ZN(n5921) );
  aoi22d1 U3911 ( .A1(n2999), .A2(n3021), .B1(memory_REGFILE_WRITE_DATA[1]), 
        .B2(n3020), .ZN(n3042) );
  aoi22d1 U3912 ( .A1(n3022), .A2(n3044), .B1(n3038), .B2(n3039), .ZN(n3745)
         );
  oai22d1 U3913 ( .A1(n6981), .A2(n3025), .B1(n314), .B2(n3023), .ZN(n3031) );
  aoi22d1 U3914 ( .A1(memory_REGFILE_WRITE_DATA[2]), .A2(n3027), .B1(n3026), 
        .B2(n3039), .ZN(n3028) );
  oaim21d1 U3915 ( .B1(n3029), .B2(memory_REGFILE_WRITE_DATA[0]), .A(n3028), 
        .ZN(n3030) );
  aoi211d1 U3916 ( .C1(n3032), .C2(n3745), .A(n3031), .B(n3030), .ZN(n3034) );
  oan211d1 U3917 ( .C1(n3036), .C2(n3035), .B(n3034), .A(n3033), .ZN(n3037) );
  aoi31d1 U3918 ( .B1(n3040), .B2(n3039), .B3(n3038), .A(n3037), .ZN(n3041) );
  oai211d1 U3919 ( .C1(n3044), .C2(n3043), .A(n3042), .B(n3041), .ZN(n5920) );
  aor21d1 U3920 ( .B1(n3238), .B2(execute_INSTRUCTION[4]), .A(n3045), .Z(n5919) );
  aoim21d1 U3921 ( .B1(n3558), .B2(execute_INSTRUCTION[3]), .A(n3046), .ZN(
        n5918) );
  aoim22d1 U3922 ( .A1(n3548), .A2(n3047), .B1(execute_INSTRUCTION[2]), .B2(
        n3558), .Z(n5917) );
  inv0d1 U3923 ( .I(n3247), .ZN(n3539) );
  aoim22d1 U3924 ( .A1(n3539), .A2(n3048), .B1(execute_INSTRUCTION[1]), .B2(
        n3558), .Z(n5916) );
  inv0d1 U3925 ( .I(n3049), .ZN(n3050) );
  inv0d0 U3926 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[31]), 
        .ZN(n3823) );
  inv0d0 U3927 ( .I(iBusWishbone_ADR[29]), .ZN(n3061) );
  aoi22d1 U3928 ( .A1(n3050), .A2(n3823), .B1(n3061), .B2(n3049), .ZN(n5915)
         );
  inv0d0 U3929 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[30]), 
        .ZN(n3821) );
  inv0d0 U3930 ( .I(iBusWishbone_ADR[28]), .ZN(n3062) );
  aoi22d1 U3931 ( .A1(n3050), .A2(n3821), .B1(n3062), .B2(n3049), .ZN(n5914)
         );
  inv0d0 U3932 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[29]), 
        .ZN(n6807) );
  inv0d0 U3933 ( .I(iBusWishbone_ADR[27]), .ZN(n3063) );
  aoi22d1 U3934 ( .A1(n3050), .A2(n6807), .B1(n3063), .B2(n3049), .ZN(n5913)
         );
  inv0d0 U3935 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[28]), 
        .ZN(n6812) );
  inv0d0 U3936 ( .I(iBusWishbone_ADR[26]), .ZN(n3064) );
  aoi22d1 U3937 ( .A1(n3050), .A2(n6812), .B1(n3064), .B2(n3049), .ZN(n5912)
         );
  inv0d0 U3938 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[27]), 
        .ZN(n6817) );
  inv0d0 U3939 ( .I(iBusWishbone_ADR[25]), .ZN(n3065) );
  aoi22d1 U3940 ( .A1(n3050), .A2(n6817), .B1(n3065), .B2(n3049), .ZN(n5911)
         );
  inv0d0 U3941 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[26]), 
        .ZN(n6822) );
  inv0d0 U3942 ( .I(iBusWishbone_ADR[24]), .ZN(n3066) );
  aoi22d1 U3943 ( .A1(n3050), .A2(n6822), .B1(n3066), .B2(n3049), .ZN(n5910)
         );
  inv0d0 U3944 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[25]), 
        .ZN(n6827) );
  inv0d0 U3945 ( .I(iBusWishbone_ADR[23]), .ZN(n3067) );
  aoi22d1 U3946 ( .A1(n3050), .A2(n6827), .B1(n3067), .B2(n3049), .ZN(n5909)
         );
  inv0d0 U3947 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[24]), 
        .ZN(n6832) );
  inv0d0 U3948 ( .I(iBusWishbone_ADR[22]), .ZN(n3068) );
  aoi22d1 U3949 ( .A1(n3050), .A2(n6832), .B1(n3068), .B2(n3049), .ZN(n5908)
         );
  inv0d0 U3950 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[23]), 
        .ZN(n6837) );
  inv0d0 U3951 ( .I(iBusWishbone_ADR[21]), .ZN(n3069) );
  aoi22d1 U3952 ( .A1(n3050), .A2(n6837), .B1(n3069), .B2(n3051), .ZN(n5907)
         );
  inv0d1 U3953 ( .I(n3049), .ZN(n3052) );
  inv0d0 U3954 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[22]), 
        .ZN(n6842) );
  inv0d0 U3955 ( .I(iBusWishbone_ADR[20]), .ZN(n3071) );
  aoi22d1 U3956 ( .A1(n3052), .A2(n6842), .B1(n3071), .B2(n3049), .ZN(n5906)
         );
  inv0d0 U3957 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[21]), 
        .ZN(n6847) );
  inv0d0 U3958 ( .I(iBusWishbone_ADR[19]), .ZN(n3072) );
  aoi22d1 U3959 ( .A1(n3052), .A2(n6847), .B1(n3072), .B2(n3049), .ZN(n5905)
         );
  inv0d0 U3960 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[20]), 
        .ZN(n6852) );
  inv0d0 U3961 ( .I(iBusWishbone_ADR[18]), .ZN(n3073) );
  aoi22d1 U3962 ( .A1(n3052), .A2(n6852), .B1(n3073), .B2(n3049), .ZN(n5904)
         );
  inv0d0 U3963 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[19]), 
        .ZN(n6857) );
  inv0d0 U3964 ( .I(iBusWishbone_ADR[17]), .ZN(n3074) );
  aoi22d1 U3965 ( .A1(n3052), .A2(n6857), .B1(n3074), .B2(n3049), .ZN(n5903)
         );
  inv0d0 U3966 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[18]), 
        .ZN(n6863) );
  inv0d0 U3967 ( .I(iBusWishbone_ADR[16]), .ZN(n3075) );
  aoi22d1 U3968 ( .A1(n3052), .A2(n6863), .B1(n3075), .B2(n3049), .ZN(n5902)
         );
  inv0d0 U3969 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[17]), 
        .ZN(n6868) );
  inv0d0 U3970 ( .I(iBusWishbone_ADR[15]), .ZN(n3076) );
  aoi22d1 U3971 ( .A1(n3052), .A2(n6868), .B1(n3076), .B2(n3049), .ZN(n5901)
         );
  inv0d0 U3972 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[16]), 
        .ZN(n6873) );
  inv0d0 U3973 ( .I(iBusWishbone_ADR[14]), .ZN(n3077) );
  aoi22d1 U3974 ( .A1(n3052), .A2(n6873), .B1(n3077), .B2(n3049), .ZN(n5900)
         );
  inv0d0 U3975 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[15]), 
        .ZN(n6880) );
  inv0d0 U3976 ( .I(iBusWishbone_ADR[13]), .ZN(n3078) );
  aoi22d1 U3977 ( .A1(n3052), .A2(n6880), .B1(n3078), .B2(n3051), .ZN(n5899)
         );
  inv0d0 U3978 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[14]), 
        .ZN(n6885) );
  inv0d0 U3979 ( .I(iBusWishbone_ADR[12]), .ZN(n3081) );
  aoi22d1 U3980 ( .A1(n3052), .A2(n6885), .B1(n3081), .B2(n3049), .ZN(n5898)
         );
  inv0d0 U3981 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[13]), 
        .ZN(n6891) );
  inv0d0 U3982 ( .I(iBusWishbone_ADR[11]), .ZN(n3082) );
  aoi22d1 U3983 ( .A1(n3052), .A2(n6891), .B1(n3082), .B2(n3049), .ZN(n5897)
         );
  inv0d0 U3984 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[12]), 
        .ZN(n3819) );
  inv0d0 U3985 ( .I(iBusWishbone_ADR[10]), .ZN(n3083) );
  aoi22d1 U3986 ( .A1(n3050), .A2(n3819), .B1(n3083), .B2(n3051), .ZN(n5896)
         );
  inv0d0 U3987 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[11]), 
        .ZN(n6898) );
  inv0d0 U3988 ( .I(iBusWishbone_ADR[9]), .ZN(n3084) );
  aoi22d1 U3989 ( .A1(n3050), .A2(n6898), .B1(n3084), .B2(n3051), .ZN(n5895)
         );
  inv0d0 U3990 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[10]), 
        .ZN(n6903) );
  inv0d0 U3991 ( .I(iBusWishbone_ADR[8]), .ZN(n3085) );
  aoi22d1 U3992 ( .A1(n3052), .A2(n6903), .B1(n3085), .B2(n3051), .ZN(n5894)
         );
  inv0d0 U3993 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[9]), 
        .ZN(n6909) );
  inv0d0 U3994 ( .I(iBusWishbone_ADR[7]), .ZN(n3086) );
  aoi22d1 U3995 ( .A1(n3050), .A2(n6909), .B1(n3086), .B2(n3051), .ZN(n5893)
         );
  inv0d0 U3996 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[8]), 
        .ZN(n6914) );
  inv0d0 U3997 ( .I(iBusWishbone_ADR[6]), .ZN(n3087) );
  aoi22d1 U3998 ( .A1(n3052), .A2(n6914), .B1(n3087), .B2(n3051), .ZN(n5892)
         );
  inv0d0 U3999 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[7]), 
        .ZN(n6924) );
  inv0d0 U4000 ( .I(iBusWishbone_ADR[5]), .ZN(n3088) );
  aoi22d1 U4001 ( .A1(n3050), .A2(n6924), .B1(n3088), .B2(n3051), .ZN(n5891)
         );
  inv0d0 U4002 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[6]), 
        .ZN(n6937) );
  inv0d0 U4003 ( .I(iBusWishbone_ADR[4]), .ZN(n3090) );
  aoi22d1 U4004 ( .A1(n3052), .A2(n6937), .B1(n3090), .B2(n3051), .ZN(n5890)
         );
  inv0d0 U4005 ( .I(IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[5]), 
        .ZN(n7000) );
  aoi22d1 U4006 ( .A1(n3052), .A2(n7000), .B1(\iBusWishbone_ADR[3]_BAR ), .B2(
        n3051), .ZN(n5889) );
  inv0d0 U4007 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][0] ), .ZN(n7010) );
  nd02d0 U4008 ( .A1(iBusWishbone_ADR[3]), .A2(n3059), .ZN(n3121) );
  nr02d0 U4009 ( .A1(n3138), .A2(n3121), .ZN(n3092) );
  buffd1 U4010 ( .I(n3092), .Z(n3093) );
  nd02d0 U4011 ( .A1(\IBusCachedPlugin_cache/_zz_ways_0_tags_port[0] ), .A2(
        n3093), .ZN(n3053) );
  aon211d1 U4012 ( .C1(\IBusCachedPlugin_cache/lineLoader_flushCounter[0] ), 
        .C2(n3054), .B(n7010), .A(n3053), .ZN(n5888) );
  buffd1 U4013 ( .I(n3092), .Z(n3096) );
  aoi22d1 U4014 ( .A1(\IBusCachedPlugin_cache/_zz_ways_0_tags_port[0] ), .A2(
        n3096), .B1(\IBusCachedPlugin_cache/lineLoader_flushCounter[0] ), .B2(
        n3054), .ZN(n3055) );
  inv0d1 U4015 ( .I(n3055), .ZN(n3057) );
  inv0d0 U4016 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][27] ), .ZN(n7011)
         );
  inv0d1 U4017 ( .I(n3055), .ZN(n3056) );
  aoi22d1 U4018 ( .A1(n3058), .A2(n7011), .B1(n3061), .B2(n3056), .ZN(n5887)
         );
  inv0d0 U4019 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][26] ), .ZN(n7014)
         );
  aoi22d1 U4020 ( .A1(n3055), .A2(n7014), .B1(n3062), .B2(n3056), .ZN(n5886)
         );
  inv0d0 U4021 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][25] ), .ZN(n7019)
         );
  aoi22d1 U4022 ( .A1(n3055), .A2(n7019), .B1(n3063), .B2(n3056), .ZN(n5885)
         );
  inv0d0 U4023 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][24] ), .ZN(n7022)
         );
  aoi22d1 U4024 ( .A1(n3055), .A2(n7022), .B1(n3064), .B2(n3056), .ZN(n5884)
         );
  inv0d0 U4025 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][23] ), .ZN(n7023)
         );
  aoi22d1 U4026 ( .A1(n3058), .A2(n7023), .B1(n3065), .B2(n3056), .ZN(n5883)
         );
  inv0d0 U4027 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][22] ), .ZN(n7028)
         );
  aoi22d1 U4028 ( .A1(n3055), .A2(n7028), .B1(n3066), .B2(n3056), .ZN(n5882)
         );
  inv0d0 U4029 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][21] ), .ZN(n7031)
         );
  aoi22d1 U4030 ( .A1(n3055), .A2(n7031), .B1(n3067), .B2(n3056), .ZN(n5881)
         );
  inv0d0 U4031 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][20] ), .ZN(n7034)
         );
  aoi22d1 U4032 ( .A1(n3055), .A2(n7034), .B1(n3068), .B2(n3056), .ZN(n5880)
         );
  inv0d0 U4033 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][19] ), .ZN(n7035)
         );
  aoi22d1 U4034 ( .A1(n3055), .A2(n7035), .B1(n3069), .B2(n3056), .ZN(n5879)
         );
  inv0d0 U4035 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][18] ), .ZN(n7040)
         );
  aoi22d1 U4036 ( .A1(n3055), .A2(n7040), .B1(n3071), .B2(n3056), .ZN(n5878)
         );
  inv0d0 U4037 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][17] ), .ZN(n7043)
         );
  aoi22d1 U4038 ( .A1(n3055), .A2(n7043), .B1(n3072), .B2(n3056), .ZN(n5877)
         );
  inv0d0 U4039 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][16] ), .ZN(n7046)
         );
  aoi22d1 U4040 ( .A1(n3055), .A2(n7046), .B1(n3073), .B2(n3056), .ZN(n5876)
         );
  inv0d0 U4041 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][15] ), .ZN(n7047)
         );
  aoi22d1 U4042 ( .A1(n3055), .A2(n7047), .B1(n3074), .B2(n3057), .ZN(n5875)
         );
  inv0d0 U4043 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][14] ), .ZN(n7052)
         );
  aoi22d1 U4044 ( .A1(n3055), .A2(n7052), .B1(n3075), .B2(n3057), .ZN(n5874)
         );
  inv0d0 U4045 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][13] ), .ZN(n7053)
         );
  aoi22d1 U4046 ( .A1(n3055), .A2(n7053), .B1(n3076), .B2(n3057), .ZN(n5873)
         );
  inv0d0 U4047 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][12] ), .ZN(n7056)
         );
  aoi22d1 U4048 ( .A1(n3055), .A2(n7056), .B1(n3077), .B2(n3057), .ZN(n5872)
         );
  inv0d0 U4049 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][11] ), .ZN(n7059)
         );
  aoi22d1 U4050 ( .A1(n3058), .A2(n7059), .B1(n3078), .B2(n3057), .ZN(n5871)
         );
  inv0d0 U4051 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][10] ), .ZN(n7064)
         );
  aoi22d1 U4052 ( .A1(n3058), .A2(n7064), .B1(n3081), .B2(n3057), .ZN(n5870)
         );
  inv0d0 U4053 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][9] ), .ZN(n7065) );
  aoi22d1 U4054 ( .A1(n3058), .A2(n7065), .B1(n3082), .B2(n3057), .ZN(n5869)
         );
  inv0d0 U4055 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][8] ), .ZN(n7068) );
  aoi22d1 U4056 ( .A1(n3058), .A2(n7068), .B1(n3083), .B2(n3057), .ZN(n5868)
         );
  inv0d0 U4057 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][7] ), .ZN(n7071) );
  aoi22d1 U4058 ( .A1(n3058), .A2(n7071), .B1(n3084), .B2(n3057), .ZN(n5867)
         );
  inv0d0 U4059 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][6] ), .ZN(n7076) );
  aoi22d1 U4060 ( .A1(n3058), .A2(n7076), .B1(n3085), .B2(n3057), .ZN(n5866)
         );
  inv0d0 U4061 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][5] ), .ZN(n7080) );
  aoi22d1 U4062 ( .A1(n3058), .A2(n7080), .B1(n3086), .B2(n3057), .ZN(n5865)
         );
  inv0d0 U4063 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][4] ), .ZN(n7083) );
  aoi22d1 U4064 ( .A1(n3058), .A2(n7083), .B1(n3087), .B2(n3057), .ZN(n5864)
         );
  inv0d0 U4065 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][3] ), .ZN(n7088) );
  aoi22d1 U4066 ( .A1(n3058), .A2(n7088), .B1(n3088), .B2(n3057), .ZN(n5863)
         );
  inv0d0 U4067 ( .I(\IBusCachedPlugin_cache/ways_0_tags[1][2] ), .ZN(n7093) );
  aoi22d1 U4068 ( .A1(n3058), .A2(n7093), .B1(n3090), .B2(n3057), .ZN(n5862)
         );
  inv0d0 U4069 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][0] ), .ZN(n7008) );
  nd02d0 U4070 ( .A1(n3059), .A2(\iBusWishbone_ADR[3]_BAR ), .ZN(n3165) );
  nr02d0 U4071 ( .A1(n3138), .A2(n3165), .ZN(n3133) );
  buffd1 U4072 ( .I(n3133), .Z(n3135) );
  oaim22d1 U4073 ( .A1(n3060), .A2(n7008), .B1(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port[0] ), .B2(n3135), .ZN(
        n5861) );
  aoi21d1 U4074 ( .B1(n3135), .B2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port[0] ), .A(n3060), .ZN(
        n3079) );
  inv0d1 U4075 ( .I(n3079), .ZN(n3089) );
  inv0d0 U4076 ( .I(n3089), .ZN(n3070) );
  inv0d0 U4077 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][27] ), .ZN(n7013)
         );
  inv0d1 U4078 ( .I(n3079), .ZN(n3080) );
  aoi22d1 U4079 ( .A1(n3070), .A2(n7013), .B1(n3061), .B2(n3080), .ZN(n5860)
         );
  inv0d0 U4080 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][26] ), .ZN(n7016)
         );
  aoi22d1 U4081 ( .A1(n3070), .A2(n7016), .B1(n3062), .B2(n3080), .ZN(n5859)
         );
  inv0d0 U4082 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][25] ), .ZN(n7017)
         );
  aoi22d1 U4083 ( .A1(n3070), .A2(n7017), .B1(n3063), .B2(n3080), .ZN(n5858)
         );
  inv0d0 U4084 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][24] ), .ZN(n7020)
         );
  aoi22d1 U4085 ( .A1(n3070), .A2(n7020), .B1(n3064), .B2(n3080), .ZN(n5857)
         );
  inv0d0 U4086 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][23] ), .ZN(n7025)
         );
  aoi22d1 U4087 ( .A1(n3070), .A2(n7025), .B1(n3065), .B2(n3080), .ZN(n5856)
         );
  inv0d0 U4088 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][22] ), .ZN(n7026)
         );
  aoi22d1 U4089 ( .A1(n3070), .A2(n7026), .B1(n3066), .B2(n3080), .ZN(n5855)
         );
  inv0d0 U4090 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][21] ), .ZN(n7029)
         );
  aoi22d1 U4091 ( .A1(n3070), .A2(n7029), .B1(n3067), .B2(n3080), .ZN(n5854)
         );
  inv0d0 U4092 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][20] ), .ZN(n7032)
         );
  aoi22d1 U4093 ( .A1(n3070), .A2(n7032), .B1(n3068), .B2(n3080), .ZN(n5853)
         );
  inv0d0 U4094 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][19] ), .ZN(n7037)
         );
  aoi22d1 U4095 ( .A1(n3070), .A2(n7037), .B1(n3069), .B2(n3080), .ZN(n5852)
         );
  inv0d0 U4096 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][18] ), .ZN(n7038)
         );
  aoi22d1 U4097 ( .A1(n3079), .A2(n7038), .B1(n3071), .B2(n3080), .ZN(n5851)
         );
  inv0d0 U4098 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][17] ), .ZN(n7041)
         );
  aoi22d1 U4099 ( .A1(n3079), .A2(n7041), .B1(n3072), .B2(n3080), .ZN(n5850)
         );
  inv0d0 U4100 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][16] ), .ZN(n7044)
         );
  aoi22d1 U4101 ( .A1(n3079), .A2(n7044), .B1(n3073), .B2(n3080), .ZN(n5849)
         );
  inv0d0 U4102 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][15] ), .ZN(n7049)
         );
  aoi22d1 U4103 ( .A1(n3079), .A2(n7049), .B1(n3074), .B2(n3089), .ZN(n5848)
         );
  inv0d0 U4104 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][14] ), .ZN(n7050)
         );
  aoi22d1 U4105 ( .A1(n3079), .A2(n7050), .B1(n3075), .B2(n3089), .ZN(n5847)
         );
  inv0d0 U4106 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][13] ), .ZN(n7055)
         );
  aoi22d1 U4107 ( .A1(n3079), .A2(n7055), .B1(n3076), .B2(n3089), .ZN(n5846)
         );
  inv0d0 U4108 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][12] ), .ZN(n7058)
         );
  aoi22d1 U4109 ( .A1(n3079), .A2(n7058), .B1(n3077), .B2(n3089), .ZN(n5845)
         );
  inv0d0 U4110 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][11] ), .ZN(n7061)
         );
  aoi22d1 U4111 ( .A1(n3079), .A2(n7061), .B1(n3078), .B2(n3089), .ZN(n5844)
         );
  inv0d0 U4112 ( .I(n3080), .ZN(n3091) );
  inv0d0 U4113 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][10] ), .ZN(n7062)
         );
  aoi22d1 U4114 ( .A1(n3091), .A2(n7062), .B1(n3081), .B2(n3089), .ZN(n5843)
         );
  inv0d0 U4115 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][9] ), .ZN(n7067) );
  aoi22d1 U4116 ( .A1(n3091), .A2(n7067), .B1(n3082), .B2(n3089), .ZN(n5842)
         );
  inv0d0 U4117 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][8] ), .ZN(n7070) );
  aoi22d1 U4118 ( .A1(n3091), .A2(n7070), .B1(n3083), .B2(n3089), .ZN(n5841)
         );
  inv0d0 U4119 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][7] ), .ZN(n7073) );
  aoi22d1 U4120 ( .A1(n3091), .A2(n7073), .B1(n3084), .B2(n3089), .ZN(n5840)
         );
  inv0d0 U4121 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][6] ), .ZN(n7074) );
  aoi22d1 U4122 ( .A1(n3091), .A2(n7074), .B1(n3085), .B2(n3089), .ZN(n5839)
         );
  inv0d0 U4123 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][5] ), .ZN(n7078) );
  aoi22d1 U4124 ( .A1(n3091), .A2(n7078), .B1(n3086), .B2(n3089), .ZN(n5838)
         );
  inv0d0 U4125 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][4] ), .ZN(n7081) );
  aoi22d1 U4126 ( .A1(n3091), .A2(n7081), .B1(n3087), .B2(n3089), .ZN(n5837)
         );
  inv0d0 U4127 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][3] ), .ZN(n7084) );
  aoi22d1 U4128 ( .A1(n3091), .A2(n7084), .B1(n3088), .B2(n3089), .ZN(n5836)
         );
  inv0d0 U4129 ( .I(\IBusCachedPlugin_cache/ways_0_tags[0][2] ), .ZN(n7089) );
  aoi22d1 U4130 ( .A1(n3091), .A2(n7089), .B1(n3090), .B2(n3089), .ZN(n5835)
         );
  inv0d1 U4131 ( .I(iBus_rsp_payload_data[0]), .ZN(n3172) );
  aoim22d1 U4132 ( .A1(n3093), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[15][0] ), .B2(n3093), .Z(n5834) );
  buffd1 U4133 ( .I(n3092), .Z(n3094) );
  aoim22d1 U4134 ( .A1(n3094), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[15][31] ), .B2(n3093), .Z(n5833) );
  buffd1 U4135 ( .I(n3092), .Z(n3095) );
  aoim22d1 U4136 ( .A1(n3095), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[15][30] ), .B2(n3093), .Z(n5832) );
  aoim22d1 U4137 ( .A1(n3094), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[15][29] ), .B2(n3093), .Z(n5831) );
  aoim22d1 U4138 ( .A1(n3093), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[15][28] ), .B2(n3093), .Z(n5830) );
  aoim22d1 U4139 ( .A1(n3095), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[15][27] ), .B2(n3093), .Z(n5829) );
  aoim22d1 U4140 ( .A1(n3094), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[15][26] ), .B2(n3093), .Z(n5828) );
  aoim22d1 U4141 ( .A1(n3093), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[15][25] ), .B2(n3095), .Z(n5827) );
  aoim22d1 U4142 ( .A1(n3095), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[15][24] ), .B2(n3093), .Z(n5826) );
  inv0d1 U4143 ( .I(iBus_rsp_payload_data[23]), .ZN(n3180) );
  aoim22d1 U4144 ( .A1(n3093), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[15][23] ), .B2(n3094), .Z(n5825) );
  inv0d1 U4145 ( .I(iBus_rsp_payload_data[22]), .ZN(n3181) );
  aoim22d1 U4146 ( .A1(n3093), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[15][22] ), .B2(n3094), .Z(n5824) );
  inv0d1 U4147 ( .I(iBus_rsp_payload_data[21]), .ZN(n3182) );
  aoim22d1 U4148 ( .A1(n3094), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[15][21] ), .B2(n3094), .Z(n5823) );
  inv0d1 U4149 ( .I(iBus_rsp_payload_data[20]), .ZN(n3183) );
  aoim22d1 U4150 ( .A1(n3093), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[15][20] ), .B2(n3094), .Z(n5822) );
  inv0d1 U4151 ( .I(iBus_rsp_payload_data[19]), .ZN(n3184) );
  aoim22d1 U4152 ( .A1(n3095), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[15][19] ), .B2(n3094), .Z(n5821) );
  inv0d1 U4153 ( .I(iBus_rsp_payload_data[18]), .ZN(n3185) );
  aoim22d1 U4154 ( .A1(n3096), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[15][18] ), .B2(n3094), .Z(n5820) );
  inv0d1 U4155 ( .I(iBus_rsp_payload_data[17]), .ZN(n3186) );
  aoim22d1 U4156 ( .A1(n3096), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[15][17] ), .B2(n3094), .Z(n5819) );
  inv0d1 U4157 ( .I(iBus_rsp_payload_data[16]), .ZN(n3187) );
  aoim22d1 U4158 ( .A1(n3096), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[15][16] ), .B2(n3094), .Z(n5818) );
  inv0d1 U4159 ( .I(iBus_rsp_payload_data[15]), .ZN(n3188) );
  aoim22d1 U4160 ( .A1(n3095), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[15][15] ), .B2(n3094), .Z(n5817) );
  inv0d1 U4161 ( .I(iBus_rsp_payload_data[14]), .ZN(n3189) );
  aoim22d1 U4162 ( .A1(n3096), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[15][14] ), .B2(n3094), .Z(n5816) );
  inv0d1 U4163 ( .I(iBus_rsp_payload_data[13]), .ZN(n3190) );
  aoim22d1 U4164 ( .A1(n3096), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[15][13] ), .B2(n3095), .Z(n5815) );
  inv0d1 U4165 ( .I(iBus_rsp_payload_data[12]), .ZN(n3193) );
  aoim22d1 U4166 ( .A1(n3093), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[15][12] ), .B2(n3095), .Z(n5814) );
  inv0d1 U4167 ( .I(iBus_rsp_payload_data[11]), .ZN(n3194) );
  aoim22d1 U4168 ( .A1(n3094), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[15][11] ), .B2(n3095), .Z(n5813) );
  inv0d1 U4169 ( .I(iBus_rsp_payload_data[10]), .ZN(n3195) );
  aoim22d1 U4170 ( .A1(n3096), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[15][10] ), .B2(n3095), .Z(n5812) );
  inv0d1 U4171 ( .I(iBus_rsp_payload_data[9]), .ZN(n3196) );
  aoim22d1 U4172 ( .A1(n3094), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[15][9] ), .B2(n3095), .Z(n5811) );
  inv0d1 U4173 ( .I(iBus_rsp_payload_data[8]), .ZN(n3198) );
  aoim22d1 U4174 ( .A1(n3095), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[15][8] ), .B2(n3095), .Z(n5810) );
  inv0d1 U4175 ( .I(iBus_rsp_payload_data[7]), .ZN(n3199) );
  aoim22d1 U4176 ( .A1(n3093), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[15][7] ), .B2(n3095), .Z(n5809) );
  inv0d1 U4177 ( .I(iBus_rsp_payload_data[6]), .ZN(n3200) );
  aoim22d1 U4178 ( .A1(n3094), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[15][6] ), .B2(n3095), .Z(n5808) );
  inv0d1 U4179 ( .I(iBus_rsp_payload_data[5]), .ZN(n3201) );
  aoim22d1 U4180 ( .A1(n3095), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[15][5] ), .B2(n3096), .Z(n5807) );
  inv0d1 U4181 ( .I(iBus_rsp_payload_data[4]), .ZN(n3202) );
  aoim22d1 U4182 ( .A1(n3096), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[15][4] ), .B2(n3096), .Z(n5806) );
  inv0d1 U4183 ( .I(iBus_rsp_payload_data[3]), .ZN(n3203) );
  aoim22d1 U4184 ( .A1(n3096), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[15][3] ), .B2(n3096), .Z(n5805) );
  inv0d1 U4185 ( .I(iBus_rsp_payload_data[2]), .ZN(n3204) );
  aoim22d1 U4186 ( .A1(n3096), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[15][2] ), .B2(n3095), .Z(n5804) );
  inv0d1 U4187 ( .I(iBus_rsp_payload_data[1]), .ZN(n3206) );
  aoim22d1 U4188 ( .A1(n3096), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[15][1] ), .B2(n3096), .Z(n5803) );
  nd03d0 U4189 ( .A1(iBusWishbone_ADR[3]), .A2(iBus_rsp_valid), .A3(n3097), 
        .ZN(n3127) );
  nr02d1 U4190 ( .A1(n3138), .A2(n3127), .ZN(n3098) );
  buffd1 U4191 ( .I(n3098), .Z(n3099) );
  buffd1 U4192 ( .I(n3098), .Z(n3101) );
  aoim22d1 U4193 ( .A1(n3099), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[14][0] ), .B2(n3101), .Z(n5802) );
  aoim22d1 U4194 ( .A1(n3100), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[14][31] ), .B2(n3101), .Z(n5801) );
  aoim22d1 U4195 ( .A1(n3099), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[14][30] ), .B2(n3101), .Z(n5800) );
  aoim22d1 U4196 ( .A1(n3099), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[14][29] ), .B2(n3098), .Z(n5799) );
  buffd1 U4197 ( .I(n3098), .Z(n3100) );
  aoim22d1 U4198 ( .A1(n3100), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[14][28] ), .B2(n3098), .Z(n5798) );
  aoim22d1 U4199 ( .A1(n3099), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[14][27] ), .B2(n3100), .Z(n5797) );
  aoim22d1 U4200 ( .A1(n3099), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[14][26] ), .B2(n3099), .Z(n5796) );
  aoim22d1 U4201 ( .A1(n3098), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[14][25] ), .B2(n3100), .Z(n5795) );
  aoim22d1 U4202 ( .A1(n3098), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[14][24] ), .B2(n3099), .Z(n5794) );
  aoim22d1 U4203 ( .A1(n3099), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[14][23] ), .B2(n3100), .Z(n5793) );
  aoim22d1 U4204 ( .A1(n3099), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[14][22] ), .B2(n3099), .Z(n5792) );
  aoim22d1 U4205 ( .A1(n3099), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[14][21] ), .B2(n3099), .Z(n5791) );
  aoim22d1 U4206 ( .A1(n3098), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[14][20] ), .B2(n3100), .Z(n5790) );
  aoim22d1 U4207 ( .A1(n3100), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[14][19] ), .B2(n3099), .Z(n5789) );
  aoim22d1 U4208 ( .A1(n3101), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[14][18] ), .B2(n3099), .Z(n5788) );
  aoim22d1 U4209 ( .A1(n3100), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[14][17] ), .B2(n3100), .Z(n5787) );
  aoim22d1 U4210 ( .A1(n3099), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[14][16] ), .B2(n3100), .Z(n5786) );
  aoim22d1 U4211 ( .A1(n3098), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[14][15] ), .B2(n3100), .Z(n5785) );
  aoim22d1 U4212 ( .A1(n3100), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[14][14] ), .B2(n3100), .Z(n5784) );
  aoim22d1 U4213 ( .A1(n3101), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[14][13] ), .B2(n3100), .Z(n5783) );
  aoim22d1 U4214 ( .A1(n3099), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[14][12] ), .B2(n3100), .Z(n5782) );
  aoim22d1 U4215 ( .A1(n3101), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[14][11] ), .B2(n3098), .Z(n5781) );
  aoim22d1 U4216 ( .A1(n3101), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[14][10] ), .B2(n3098), .Z(n5780) );
  aoim22d1 U4217 ( .A1(n3098), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[14][9] ), .B2(n3098), .Z(n5779) );
  aoim22d1 U4218 ( .A1(n3101), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[14][8] ), .B2(n3098), .Z(n5778) );
  aoim22d1 U4219 ( .A1(n3100), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[14][7] ), .B2(n3098), .Z(n5777) );
  aoim22d1 U4220 ( .A1(n3101), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[14][6] ), .B2(n3098), .Z(n5776) );
  aoim22d1 U4221 ( .A1(n3101), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[14][5] ), .B2(n3101), .Z(n5775) );
  aoim22d1 U4222 ( .A1(n3099), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[14][4] ), .B2(n3101), .Z(n5774) );
  aoim22d1 U4223 ( .A1(n3100), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[14][3] ), .B2(n3101), .Z(n5773) );
  aoim22d1 U4224 ( .A1(n3101), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[14][2] ), .B2(n3101), .Z(n5772) );
  aoim22d1 U4225 ( .A1(n3101), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[14][1] ), .B2(n3101), .Z(n5771) );
  buffd1 U4226 ( .I(n3102), .Z(n3104) );
  buffd1 U4227 ( .I(n3102), .Z(n3106) );
  aoim22d1 U4228 ( .A1(n3104), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[13][0] ), .B2(n3106), .Z(n5770) );
  buffd1 U4229 ( .I(n3102), .Z(n3103) );
  aoim22d1 U4230 ( .A1(n3103), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[13][31] ), .B2(n3106), .Z(n5769) );
  aoim22d1 U4231 ( .A1(n3104), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[13][30] ), .B2(n3103), .Z(n5768) );
  aoim22d1 U4232 ( .A1(n3104), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[13][29] ), .B2(n3103), .Z(n5767) );
  buffd1 U4233 ( .I(n3102), .Z(n3105) );
  aoim22d1 U4234 ( .A1(n3105), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[13][28] ), .B2(n3103), .Z(n5766) );
  aoim22d1 U4235 ( .A1(n3104), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[13][27] ), .B2(n3105), .Z(n5765) );
  aoim22d1 U4236 ( .A1(n3104), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[13][26] ), .B2(n3103), .Z(n5764) );
  aoim22d1 U4237 ( .A1(n3103), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[13][25] ), .B2(n3105), .Z(n5763) );
  aoim22d1 U4238 ( .A1(n3103), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[13][24] ), .B2(n3104), .Z(n5762) );
  aoim22d1 U4239 ( .A1(n3104), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[13][23] ), .B2(n3105), .Z(n5761) );
  aoim22d1 U4240 ( .A1(n3104), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[13][22] ), .B2(n3104), .Z(n5760) );
  aoim22d1 U4241 ( .A1(n3104), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[13][21] ), .B2(n3104), .Z(n5759) );
  aoim22d1 U4242 ( .A1(n3103), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[13][20] ), .B2(n3105), .Z(n5758) );
  aoim22d1 U4243 ( .A1(n3105), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[13][19] ), .B2(n3104), .Z(n5757) );
  aoim22d1 U4244 ( .A1(n3106), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[13][18] ), .B2(n3104), .Z(n5756) );
  aoim22d1 U4245 ( .A1(n3105), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[13][17] ), .B2(n3105), .Z(n5755) );
  aoim22d1 U4246 ( .A1(n3104), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[13][16] ), .B2(n3105), .Z(n5754) );
  aoim22d1 U4247 ( .A1(n3103), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[13][15] ), .B2(n3105), .Z(n5753) );
  aoim22d1 U4248 ( .A1(n3105), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[13][14] ), .B2(n3105), .Z(n5752) );
  aoim22d1 U4249 ( .A1(n3106), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[13][13] ), .B2(n3105), .Z(n5751) );
  aoim22d1 U4250 ( .A1(n3104), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[13][12] ), .B2(n3105), .Z(n5750) );
  aoim22d1 U4251 ( .A1(n3106), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[13][11] ), .B2(n3103), .Z(n5749) );
  aoim22d1 U4252 ( .A1(n3106), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[13][10] ), .B2(n3103), .Z(n5748) );
  aoim22d1 U4253 ( .A1(n3103), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[13][9] ), .B2(n3103), .Z(n5747) );
  aoim22d1 U4254 ( .A1(n3106), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[13][8] ), .B2(n3103), .Z(n5746) );
  aoim22d1 U4255 ( .A1(n3105), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[13][7] ), .B2(n3103), .Z(n5745) );
  aoim22d1 U4256 ( .A1(n3106), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[13][6] ), .B2(n3103), .Z(n5744) );
  aoim22d1 U4257 ( .A1(n3106), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[13][5] ), .B2(n3106), .Z(n5743) );
  aoim22d1 U4258 ( .A1(n3104), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[13][4] ), .B2(n3106), .Z(n5742) );
  aoim22d1 U4259 ( .A1(n3105), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[13][3] ), .B2(n3106), .Z(n5741) );
  aoim22d1 U4260 ( .A1(n3106), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[13][2] ), .B2(n3106), .Z(n5740) );
  aoim22d1 U4261 ( .A1(n3106), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[13][1] ), .B2(n3106), .Z(n5739) );
  nr02d1 U4262 ( .A1(n3127), .A2(n3147), .ZN(n3107) );
  buffd1 U4263 ( .I(n3107), .Z(n3109) );
  buffd1 U4264 ( .I(n3107), .Z(n3110) );
  aoim22d1 U4265 ( .A1(n3109), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[12][0] ), .B2(n3110), .Z(n5738) );
  buffd1 U4266 ( .I(n3107), .Z(n3108) );
  aoim22d1 U4267 ( .A1(n3108), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[12][31] ), .B2(n3110), .Z(n5737) );
  aoim22d1 U4268 ( .A1(n3109), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[12][30] ), .B2(n3108), .Z(n5736) );
  aoim22d1 U4269 ( .A1(n3109), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[12][29] ), .B2(n3108), .Z(n5735) );
  aoim22d1 U4270 ( .A1(n3107), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[12][28] ), .B2(n3108), .Z(n5734) );
  aoim22d1 U4271 ( .A1(n3109), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[12][27] ), .B2(n3107), .Z(n5733) );
  aoim22d1 U4272 ( .A1(n3109), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[12][26] ), .B2(n3108), .Z(n5732) );
  aoim22d1 U4273 ( .A1(n3108), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[12][25] ), .B2(n3107), .Z(n5731) );
  aoim22d1 U4274 ( .A1(n3108), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[12][24] ), .B2(n3109), .Z(n5730) );
  aoim22d1 U4275 ( .A1(n3109), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[12][23] ), .B2(n3107), .Z(n5729) );
  aoim22d1 U4276 ( .A1(n3109), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[12][22] ), .B2(n3109), .Z(n5728) );
  aoim22d1 U4277 ( .A1(n3109), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[12][21] ), .B2(n3109), .Z(n5727) );
  aoim22d1 U4278 ( .A1(n3108), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[12][20] ), .B2(n3107), .Z(n5726) );
  aoim22d1 U4279 ( .A1(n3107), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[12][19] ), .B2(n3109), .Z(n5725) );
  aoim22d1 U4280 ( .A1(n3110), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[12][18] ), .B2(n3109), .Z(n5724) );
  aoim22d1 U4281 ( .A1(n3107), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[12][17] ), .B2(n3107), .Z(n5723) );
  aoim22d1 U4282 ( .A1(n3109), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[12][16] ), .B2(n3108), .Z(n5722) );
  aoim22d1 U4283 ( .A1(n3108), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[12][15] ), .B2(n3109), .Z(n5721) );
  aoim22d1 U4284 ( .A1(n3107), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[12][14] ), .B2(n3107), .Z(n5720) );
  aoim22d1 U4285 ( .A1(n3110), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[12][13] ), .B2(n3107), .Z(n5719) );
  aoim22d1 U4286 ( .A1(n3109), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[12][12] ), .B2(n3107), .Z(n5718) );
  aoim22d1 U4287 ( .A1(n3110), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[12][11] ), .B2(n3108), .Z(n5717) );
  aoim22d1 U4288 ( .A1(n3110), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[12][10] ), .B2(n3108), .Z(n5716) );
  aoim22d1 U4289 ( .A1(n3108), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[12][9] ), .B2(n3108), .Z(n5715) );
  aoim22d1 U4290 ( .A1(n3110), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[12][8] ), .B2(n3108), .Z(n5714) );
  aoim22d1 U4291 ( .A1(n3110), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[12][7] ), .B2(n3108), .Z(n5713) );
  aoim22d1 U4292 ( .A1(n3110), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[12][6] ), .B2(n3108), .Z(n5712) );
  aoim22d1 U4293 ( .A1(n3110), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[12][5] ), .B2(n3110), .Z(n5711) );
  aoim22d1 U4294 ( .A1(n3109), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[12][4] ), .B2(n3110), .Z(n5710) );
  aoim22d1 U4295 ( .A1(n3107), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[12][3] ), .B2(n3110), .Z(n5709) );
  aoim22d1 U4296 ( .A1(n3110), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[12][2] ), .B2(n3110), .Z(n5708) );
  aoim22d1 U4297 ( .A1(n3110), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[12][1] ), .B2(n3110), .Z(n5707) );
  nr03d0 U4298 ( .A1(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[2] ), 
        .A2(n3159), .A3(n3121), .ZN(n3111) );
  buffd1 U4299 ( .I(n3111), .Z(n3114) );
  buffd1 U4300 ( .I(n3111), .Z(n3113) );
  aoim22d1 U4301 ( .A1(n3114), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[11][0] ), .B2(n3113), .Z(n5706) );
  buffd1 U4302 ( .I(n3111), .Z(n3115) );
  buffd1 U4303 ( .I(n3111), .Z(n3112) );
  aoim22d1 U4304 ( .A1(n3115), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[11][31] ), .B2(n3112), .Z(n5705) );
  aoim22d1 U4305 ( .A1(n3114), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[11][30] ), .B2(n3112), .Z(n5704) );
  aoim22d1 U4306 ( .A1(n3114), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[11][29] ), .B2(n3112), .Z(n5703) );
  aoim22d1 U4307 ( .A1(n3113), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[11][28] ), .B2(n3112), .Z(n5702) );
  aoim22d1 U4308 ( .A1(n3114), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[11][27] ), .B2(n3113), .Z(n5701) );
  aoim22d1 U4309 ( .A1(n3114), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[11][26] ), .B2(n3112), .Z(n5700) );
  aoim22d1 U4310 ( .A1(n3114), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[11][25] ), .B2(n3113), .Z(n5699) );
  aoim22d1 U4311 ( .A1(n3115), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[11][24] ), .B2(n3114), .Z(n5698) );
  aoim22d1 U4312 ( .A1(n3114), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[11][23] ), .B2(n3113), .Z(n5697) );
  aoim22d1 U4313 ( .A1(n3115), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[11][22] ), .B2(n3114), .Z(n5696) );
  aoim22d1 U4314 ( .A1(n3115), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[11][21] ), .B2(n3114), .Z(n5695) );
  aoim22d1 U4315 ( .A1(n3112), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[11][20] ), .B2(n3113), .Z(n5694) );
  aoim22d1 U4316 ( .A1(n3115), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[11][19] ), .B2(n3114), .Z(n5693) );
  aoim22d1 U4317 ( .A1(n3115), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[11][18] ), .B2(n3114), .Z(n5692) );
  aoim22d1 U4318 ( .A1(n3113), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[11][17] ), .B2(n3113), .Z(n5691) );
  aoim22d1 U4319 ( .A1(n3115), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[11][16] ), .B2(n3113), .Z(n5690) );
  aoim22d1 U4320 ( .A1(n3115), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[11][15] ), .B2(n3113), .Z(n5689) );
  aoim22d1 U4321 ( .A1(n3115), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[11][14] ), .B2(n3113), .Z(n5688) );
  aoim22d1 U4322 ( .A1(n3115), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[11][13] ), .B2(n3113), .Z(n5687) );
  aoim22d1 U4323 ( .A1(n3115), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[11][12] ), .B2(n3113), .Z(n5686) );
  aoim22d1 U4324 ( .A1(n3115), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[11][11] ), .B2(n3112), .Z(n5685) );
  aoim22d1 U4325 ( .A1(n3115), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[11][10] ), .B2(n3112), .Z(n5684) );
  aoim22d1 U4326 ( .A1(n3115), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[11][9] ), .B2(n3112), .Z(n5683) );
  aoim22d1 U4327 ( .A1(n3112), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[11][8] ), .B2(n3112), .Z(n5682) );
  aoim22d1 U4328 ( .A1(n3112), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[11][7] ), .B2(n3112), .Z(n5681) );
  aoim22d1 U4329 ( .A1(n3112), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[11][6] ), .B2(n3112), .Z(n5680) );
  aoim22d1 U4330 ( .A1(n3112), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[11][5] ), .B2(n3114), .Z(n5679) );
  aoim22d1 U4331 ( .A1(n3113), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[11][4] ), .B2(n3113), .Z(n5678) );
  aoim22d1 U4332 ( .A1(n3114), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[11][3] ), .B2(n3114), .Z(n5677) );
  aoim22d1 U4333 ( .A1(n3115), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[11][2] ), .B2(n3113), .Z(n5676) );
  aoim22d1 U4334 ( .A1(n3115), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[11][1] ), .B2(n3114), .Z(n5675) );
  nr03d0 U4335 ( .A1(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[2] ), 
        .A2(n3159), .A3(n3127), .ZN(n3116) );
  buffd1 U4336 ( .I(n3116), .Z(n3120) );
  buffd1 U4337 ( .I(n3116), .Z(n3119) );
  aoim22d1 U4338 ( .A1(n3120), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[10][0] ), .B2(n3119), .Z(n5674) );
  buffd1 U4339 ( .I(n3116), .Z(n3117) );
  buffd1 U4340 ( .I(n3117), .Z(n3118) );
  aoim22d1 U4341 ( .A1(n3118), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[10][31] ), .B2(n3120), .Z(n5673) );
  aoim22d1 U4342 ( .A1(n3120), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[10][30] ), .B2(n3117), .Z(n5672) );
  aoim22d1 U4343 ( .A1(n3120), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[10][29] ), .B2(n3117), .Z(n5671) );
  aoim22d1 U4344 ( .A1(n3118), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[10][28] ), .B2(n3117), .Z(n5670) );
  aoim22d1 U4345 ( .A1(n3120), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[10][27] ), .B2(n3119), .Z(n5669) );
  aoim22d1 U4346 ( .A1(n3120), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[10][26] ), .B2(n3117), .Z(n5668) );
  aoim22d1 U4347 ( .A1(n3118), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[10][25] ), .B2(n3119), .Z(n5667) );
  aoim22d1 U4348 ( .A1(n3118), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[10][24] ), .B2(n3120), .Z(n5666) );
  aoim22d1 U4349 ( .A1(n3118), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[10][23] ), .B2(n3119), .Z(n5665) );
  aoim22d1 U4350 ( .A1(n3118), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[10][22] ), .B2(n3120), .Z(n5664) );
  aoim22d1 U4351 ( .A1(n3118), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[10][21] ), .B2(n3120), .Z(n5663) );
  aoim22d1 U4352 ( .A1(n3118), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[10][20] ), .B2(n3119), .Z(n5662) );
  aoim22d1 U4353 ( .A1(n3119), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[10][19] ), .B2(n3120), .Z(n5661) );
  aoim22d1 U4354 ( .A1(n3117), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[10][18] ), .B2(n3120), .Z(n5660) );
  aoim22d1 U4355 ( .A1(n3118), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[10][17] ), .B2(n3119), .Z(n5659) );
  aoim22d1 U4356 ( .A1(n3120), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[10][16] ), .B2(n3119), .Z(n5658) );
  aoim22d1 U4357 ( .A1(n3117), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[10][15] ), .B2(n3119), .Z(n5657) );
  aoim22d1 U4358 ( .A1(n3118), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[10][14] ), .B2(n3119), .Z(n5656) );
  aoim22d1 U4359 ( .A1(n3117), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[10][13] ), .B2(n3119), .Z(n5655) );
  aoim22d1 U4360 ( .A1(n3118), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[10][12] ), .B2(n3119), .Z(n5654) );
  aoim22d1 U4361 ( .A1(n3118), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[10][11] ), .B2(n3117), .Z(n5653) );
  aoim22d1 U4362 ( .A1(n3117), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[10][10] ), .B2(n3117), .Z(n5652) );
  aoim22d1 U4363 ( .A1(n3118), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[10][9] ), .B2(n3117), .Z(n5651) );
  aoim22d1 U4364 ( .A1(n3119), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[10][8] ), .B2(n3117), .Z(n5650) );
  aoim22d1 U4365 ( .A1(n3120), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[10][7] ), .B2(n3117), .Z(n5649) );
  aoim22d1 U4366 ( .A1(n3117), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[10][6] ), .B2(n3117), .Z(n5648) );
  aoim22d1 U4367 ( .A1(n3117), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[10][5] ), .B2(n3120), .Z(n5647) );
  aoim22d1 U4368 ( .A1(n3119), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[10][4] ), .B2(n3119), .Z(n5646) );
  aoim22d1 U4369 ( .A1(n3120), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[10][3] ), .B2(n3119), .Z(n5645) );
  aoim22d1 U4370 ( .A1(n3118), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[10][2] ), .B2(n3120), .Z(n5644) );
  aoim22d1 U4371 ( .A1(n3120), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[10][1] ), .B2(n3119), .Z(n5643) );
  nr03d0 U4372 ( .A1(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[1] ), 
        .A2(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[2] ), 
        .A3(n3121), .ZN(n3122) );
  buffd1 U4373 ( .I(n3122), .Z(n3126) );
  buffd1 U4374 ( .I(n3122), .Z(n3125) );
  aoim22d1 U4375 ( .A1(n3126), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[9][0] ), .B2(n3125), .Z(n5642) );
  buffd1 U4376 ( .I(n3122), .Z(n3123) );
  buffd1 U4377 ( .I(n3123), .Z(n3124) );
  aoim22d1 U4378 ( .A1(n3124), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[9][31] ), .B2(n3126), .Z(n5641) );
  aoim22d1 U4379 ( .A1(n3126), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[9][30] ), .B2(n3123), .Z(n5640) );
  aoim22d1 U4380 ( .A1(n3126), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[9][29] ), .B2(n3123), .Z(n5639) );
  aoim22d1 U4381 ( .A1(n3124), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[9][28] ), .B2(n3123), .Z(n5638) );
  aoim22d1 U4382 ( .A1(n3126), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[9][27] ), .B2(n3125), .Z(n5637) );
  aoim22d1 U4383 ( .A1(n3126), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[9][26] ), .B2(n3123), .Z(n5636) );
  aoim22d1 U4384 ( .A1(n3124), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[9][25] ), .B2(n3125), .Z(n5635) );
  aoim22d1 U4385 ( .A1(n3124), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[9][24] ), .B2(n3126), .Z(n5634) );
  aoim22d1 U4386 ( .A1(n3124), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[9][23] ), .B2(n3125), .Z(n5633) );
  aoim22d1 U4387 ( .A1(n3124), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[9][22] ), .B2(n3126), .Z(n5632) );
  aoim22d1 U4388 ( .A1(n3124), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[9][21] ), .B2(n3126), .Z(n5631) );
  aoim22d1 U4389 ( .A1(n3124), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[9][20] ), .B2(n3125), .Z(n5630) );
  aoim22d1 U4390 ( .A1(n3125), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[9][19] ), .B2(n3126), .Z(n5629) );
  aoim22d1 U4391 ( .A1(n3123), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[9][18] ), .B2(n3126), .Z(n5628) );
  aoim22d1 U4392 ( .A1(n3124), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[9][17] ), .B2(n3125), .Z(n5627) );
  aoim22d1 U4393 ( .A1(n3126), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[9][16] ), .B2(n3125), .Z(n5626) );
  aoim22d1 U4394 ( .A1(n3123), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[9][15] ), .B2(n3125), .Z(n5625) );
  aoim22d1 U4395 ( .A1(n3124), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[9][14] ), .B2(n3125), .Z(n5624) );
  aoim22d1 U4396 ( .A1(n3123), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[9][13] ), .B2(n3125), .Z(n5623) );
  aoim22d1 U4397 ( .A1(n3124), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[9][12] ), .B2(n3125), .Z(n5622) );
  aoim22d1 U4398 ( .A1(n3124), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[9][11] ), .B2(n3123), .Z(n5621) );
  aoim22d1 U4399 ( .A1(n3123), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[9][10] ), .B2(n3123), .Z(n5620) );
  aoim22d1 U4400 ( .A1(n3124), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[9][9] ), .B2(n3123), .Z(n5619) );
  aoim22d1 U4401 ( .A1(n3125), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[9][8] ), .B2(n3123), .Z(n5618) );
  aoim22d1 U4402 ( .A1(n3126), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[9][7] ), .B2(n3123), .Z(n5617) );
  aoim22d1 U4403 ( .A1(n3123), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[9][6] ), .B2(n3123), .Z(n5616) );
  aoim22d1 U4404 ( .A1(n3123), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[9][5] ), .B2(n3126), .Z(n5615) );
  aoim22d1 U4405 ( .A1(n3125), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[9][4] ), .B2(n3125), .Z(n5614) );
  aoim22d1 U4406 ( .A1(n3126), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[9][3] ), .B2(n3125), .Z(n5613) );
  aoim22d1 U4407 ( .A1(n3124), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[9][2] ), .B2(n3126), .Z(n5612) );
  aoim22d1 U4408 ( .A1(n3126), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[9][1] ), .B2(n3125), .Z(n5611) );
  nr03d0 U4409 ( .A1(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[1] ), 
        .A2(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[2] ), 
        .A3(n3127), .ZN(n3128) );
  buffd1 U4410 ( .I(n3128), .Z(n3131) );
  buffd1 U4411 ( .I(n3128), .Z(n3130) );
  aoim22d1 U4412 ( .A1(n3131), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[8][0] ), .B2(n3130), .Z(n5610) );
  buffd1 U4413 ( .I(n3128), .Z(n3132) );
  buffd1 U4414 ( .I(n3128), .Z(n3129) );
  aoim22d1 U4415 ( .A1(n3132), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[8][31] ), .B2(n3129), .Z(n5609) );
  aoim22d1 U4416 ( .A1(n3131), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[8][30] ), .B2(n3129), .Z(n5608) );
  aoim22d1 U4417 ( .A1(n3131), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[8][29] ), .B2(n3129), .Z(n5607) );
  aoim22d1 U4418 ( .A1(n3130), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[8][28] ), .B2(n3129), .Z(n5606) );
  aoim22d1 U4419 ( .A1(n3131), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[8][27] ), .B2(n3130), .Z(n5605) );
  aoim22d1 U4420 ( .A1(n3131), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[8][26] ), .B2(n3129), .Z(n5604) );
  aoim22d1 U4421 ( .A1(n3131), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[8][25] ), .B2(n3130), .Z(n5603) );
  aoim22d1 U4422 ( .A1(n3132), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[8][24] ), .B2(n3131), .Z(n5602) );
  aoim22d1 U4423 ( .A1(n3131), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[8][23] ), .B2(n3130), .Z(n5601) );
  aoim22d1 U4424 ( .A1(n3132), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[8][22] ), .B2(n3131), .Z(n5600) );
  aoim22d1 U4425 ( .A1(n3132), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[8][21] ), .B2(n3131), .Z(n5599) );
  aoim22d1 U4426 ( .A1(n3129), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[8][20] ), .B2(n3130), .Z(n5598) );
  aoim22d1 U4427 ( .A1(n3132), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[8][19] ), .B2(n3131), .Z(n5597) );
  aoim22d1 U4428 ( .A1(n3132), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[8][18] ), .B2(n3131), .Z(n5596) );
  aoim22d1 U4429 ( .A1(n3130), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[8][17] ), .B2(n3130), .Z(n5595) );
  aoim22d1 U4430 ( .A1(n3132), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[8][16] ), .B2(n3130), .Z(n5594) );
  aoim22d1 U4431 ( .A1(n3132), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[8][15] ), .B2(n3130), .Z(n5593) );
  aoim22d1 U4432 ( .A1(n3132), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[8][14] ), .B2(n3130), .Z(n5592) );
  aoim22d1 U4433 ( .A1(n3132), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[8][13] ), .B2(n3130), .Z(n5591) );
  aoim22d1 U4434 ( .A1(n3132), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[8][12] ), .B2(n3130), .Z(n5590) );
  aoim22d1 U4435 ( .A1(n3132), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[8][11] ), .B2(n3129), .Z(n5589) );
  aoim22d1 U4436 ( .A1(n3132), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[8][10] ), .B2(n3129), .Z(n5588) );
  aoim22d1 U4437 ( .A1(n3132), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[8][9] ), .B2(n3129), .Z(n5587) );
  aoim22d1 U4438 ( .A1(n3129), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[8][8] ), .B2(n3129), .Z(n5586) );
  aoim22d1 U4439 ( .A1(n3129), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[8][7] ), .B2(n3129), .Z(n5585) );
  aoim22d1 U4440 ( .A1(n3129), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[8][6] ), .B2(n3129), .Z(n5584) );
  aoim22d1 U4441 ( .A1(n3129), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[8][5] ), .B2(n3131), .Z(n5583) );
  aoim22d1 U4442 ( .A1(n3130), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[8][4] ), .B2(n3130), .Z(n5582) );
  aoim22d1 U4443 ( .A1(n3131), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[8][3] ), .B2(n3131), .Z(n5581) );
  aoim22d1 U4444 ( .A1(n3132), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[8][2] ), .B2(n3130), .Z(n5580) );
  aoim22d1 U4445 ( .A1(n3132), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[8][1] ), .B2(n3131), .Z(n5579) );
  buffd1 U4446 ( .I(n3133), .Z(n3137) );
  aoim22d1 U4447 ( .A1(n3137), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[7][0] ), .B2(n3135), .Z(n5578) );
  buffd1 U4448 ( .I(n3133), .Z(n3134) );
  aoim22d1 U4449 ( .A1(n3137), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[7][31] ), .B2(n3134), .Z(n5577) );
  buffd1 U4450 ( .I(n3133), .Z(n3136) );
  aoim22d1 U4451 ( .A1(n3136), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[7][30] ), .B2(n3134), .Z(n5576) );
  aoim22d1 U4452 ( .A1(n3137), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[7][29] ), .B2(n3134), .Z(n5575) );
  aoim22d1 U4453 ( .A1(n3136), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[7][28] ), .B2(n3134), .Z(n5574) );
  aoim22d1 U4454 ( .A1(n3134), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[7][27] ), .B2(n3134), .Z(n5573) );
  aoim22d1 U4455 ( .A1(n3137), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[7][26] ), .B2(n3134), .Z(n5572) );
  aoim22d1 U4456 ( .A1(n3137), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[7][25] ), .B2(n3136), .Z(n5571) );
  aoim22d1 U4457 ( .A1(n3134), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[7][24] ), .B2(n3134), .Z(n5570) );
  aoim22d1 U4458 ( .A1(n3134), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[7][23] ), .B2(n3134), .Z(n5569) );
  aoim22d1 U4459 ( .A1(n3134), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[7][22] ), .B2(n3134), .Z(n5568) );
  aoim22d1 U4460 ( .A1(n3135), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[7][21] ), .B2(n3137), .Z(n5567) );
  aoim22d1 U4461 ( .A1(n3135), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[7][20] ), .B2(n3137), .Z(n5566) );
  aoim22d1 U4462 ( .A1(n3135), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[7][19] ), .B2(n3137), .Z(n5565) );
  aoim22d1 U4463 ( .A1(n3134), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[7][18] ), .B2(n3137), .Z(n5564) );
  aoim22d1 U4464 ( .A1(n3135), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[7][17] ), .B2(n3137), .Z(n5563) );
  aoim22d1 U4465 ( .A1(n3134), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[7][16] ), .B2(n3137), .Z(n5562) );
  aoim22d1 U4466 ( .A1(n3135), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[7][15] ), .B2(n3137), .Z(n5561) );
  aoim22d1 U4467 ( .A1(n3135), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[7][14] ), .B2(n3137), .Z(n5560) );
  aoim22d1 U4468 ( .A1(n3135), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[7][13] ), .B2(n3137), .Z(n5559) );
  aoim22d1 U4469 ( .A1(n3135), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[7][12] ), .B2(n3137), .Z(n5558) );
  aoim22d1 U4470 ( .A1(n3134), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[7][11] ), .B2(n3136), .Z(n5557) );
  aoim22d1 U4471 ( .A1(n3134), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[7][10] ), .B2(n3136), .Z(n5556) );
  aoim22d1 U4472 ( .A1(n3135), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[7][9] ), .B2(n3136), .Z(n5555) );
  aoim22d1 U4473 ( .A1(n3135), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[7][8] ), .B2(n3136), .Z(n5554) );
  aoim22d1 U4474 ( .A1(n3136), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[7][7] ), .B2(n3136), .Z(n5553) );
  aoim22d1 U4475 ( .A1(n3136), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[7][6] ), .B2(n3136), .Z(n5552) );
  aoim22d1 U4476 ( .A1(n3136), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[7][5] ), .B2(n3135), .Z(n5551) );
  aoim22d1 U4477 ( .A1(n3137), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[7][4] ), .B2(n3135), .Z(n5550) );
  aoim22d1 U4478 ( .A1(n3136), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[7][3] ), .B2(n3136), .Z(n5549) );
  aoim22d1 U4479 ( .A1(n3136), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[7][2] ), .B2(n3136), .Z(n5548) );
  aoim22d1 U4480 ( .A1(n3137), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[7][1] ), .B2(n3136), .Z(n5547) );
  nr02d1 U4481 ( .A1(n3138), .A2(n3158), .ZN(n3139) );
  buffd1 U4482 ( .I(n3139), .Z(n3142) );
  aoim22d1 U4483 ( .A1(n3139), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[6][0] ), .B2(n3142), .Z(n5546) );
  aoim22d1 U4484 ( .A1(n3142), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[6][31] ), .B2(n3142), .Z(n5545) );
  buffd1 U4485 ( .I(n3139), .Z(n3141) );
  aoim22d1 U4486 ( .A1(n3139), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[6][30] ), .B2(n3141), .Z(n5544) );
  aoim22d1 U4487 ( .A1(n3139), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[6][29] ), .B2(n3141), .Z(n5543) );
  aoim22d1 U4488 ( .A1(n3141), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[6][28] ), .B2(n3141), .Z(n5542) );
  buffd1 U4489 ( .I(n3139), .Z(n3140) );
  aoim22d1 U4490 ( .A1(n3139), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[6][27] ), .B2(n3140), .Z(n5541) );
  aoim22d1 U4491 ( .A1(n3139), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[6][26] ), .B2(n3141), .Z(n5540) );
  aoim22d1 U4492 ( .A1(n3142), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[6][25] ), .B2(n3140), .Z(n5539) );
  aoim22d1 U4493 ( .A1(n3139), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[6][24] ), .B2(n3139), .Z(n5538) );
  aoim22d1 U4494 ( .A1(n3140), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[6][23] ), .B2(n3140), .Z(n5537) );
  aoim22d1 U4495 ( .A1(n3139), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[6][22] ), .B2(n3139), .Z(n5536) );
  aoim22d1 U4496 ( .A1(n3142), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[6][21] ), .B2(n3139), .Z(n5535) );
  aoim22d1 U4497 ( .A1(n3139), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[6][20] ), .B2(n3140), .Z(n5534) );
  aoim22d1 U4498 ( .A1(n3142), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[6][19] ), .B2(n3139), .Z(n5533) );
  aoim22d1 U4499 ( .A1(n3142), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[6][18] ), .B2(n3139), .Z(n5532) );
  aoim22d1 U4500 ( .A1(n3142), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[6][17] ), .B2(n3140), .Z(n5531) );
  aoim22d1 U4501 ( .A1(n3140), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[6][16] ), .B2(n3140), .Z(n5530) );
  aoim22d1 U4502 ( .A1(n3142), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[6][15] ), .B2(n3140), .Z(n5529) );
  aoim22d1 U4503 ( .A1(n3141), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[6][14] ), .B2(n3140), .Z(n5528) );
  aoim22d1 U4504 ( .A1(n3141), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[6][13] ), .B2(n3140), .Z(n5527) );
  aoim22d1 U4505 ( .A1(n3140), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[6][12] ), .B2(n3140), .Z(n5526) );
  aoim22d1 U4506 ( .A1(n3142), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[6][11] ), .B2(n3141), .Z(n5525) );
  aoim22d1 U4507 ( .A1(n3140), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[6][10] ), .B2(n3141), .Z(n5524) );
  aoim22d1 U4508 ( .A1(n3141), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[6][9] ), .B2(n3141), .Z(n5523) );
  aoim22d1 U4509 ( .A1(n3140), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[6][8] ), .B2(n3141), .Z(n5522) );
  aoim22d1 U4510 ( .A1(n3142), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[6][7] ), .B2(n3141), .Z(n5521) );
  aoim22d1 U4511 ( .A1(n3141), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[6][6] ), .B2(n3141), .Z(n5520) );
  aoim22d1 U4512 ( .A1(n3140), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[6][5] ), .B2(n3142), .Z(n5519) );
  aoim22d1 U4513 ( .A1(n3141), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[6][4] ), .B2(n3142), .Z(n5518) );
  aoim22d1 U4514 ( .A1(n3140), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[6][3] ), .B2(n3142), .Z(n5517) );
  aoim22d1 U4515 ( .A1(n3141), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[6][2] ), .B2(n3142), .Z(n5516) );
  aoim22d1 U4516 ( .A1(n3142), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[6][1] ), .B2(n3142), .Z(n5515) );
  nr02d1 U4517 ( .A1(n3165), .A2(n3147), .ZN(n3143) );
  buffd1 U4518 ( .I(n3143), .Z(n3144) );
  buffd1 U4519 ( .I(n3143), .Z(n3146) );
  aoim22d1 U4520 ( .A1(n3144), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[5][0] ), .B2(n3146), .Z(n5514) );
  aoim22d1 U4521 ( .A1(n3146), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[5][31] ), .B2(n3146), .Z(n5513) );
  buffd1 U4522 ( .I(n3143), .Z(n3145) );
  aoim22d1 U4523 ( .A1(n3144), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[5][30] ), .B2(n3145), .Z(n5512) );
  aoim22d1 U4524 ( .A1(n3144), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[5][29] ), .B2(n3145), .Z(n5511) );
  aoim22d1 U4525 ( .A1(n3145), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[5][28] ), .B2(n3145), .Z(n5510) );
  aoim22d1 U4526 ( .A1(n3144), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[5][27] ), .B2(n3143), .Z(n5509) );
  aoim22d1 U4527 ( .A1(n3144), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[5][26] ), .B2(n3145), .Z(n5508) );
  aoim22d1 U4528 ( .A1(n3146), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[5][25] ), .B2(n3144), .Z(n5507) );
  aoim22d1 U4529 ( .A1(n3144), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[5][24] ), .B2(n3144), .Z(n5506) );
  aoim22d1 U4530 ( .A1(n3143), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[5][23] ), .B2(n3146), .Z(n5505) );
  aoim22d1 U4531 ( .A1(n3144), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[5][22] ), .B2(n3144), .Z(n5504) );
  aoim22d1 U4532 ( .A1(n3146), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[5][21] ), .B2(n3144), .Z(n5503) );
  aoim22d1 U4533 ( .A1(n3144), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[5][20] ), .B2(n3145), .Z(n5502) );
  aoim22d1 U4534 ( .A1(n3146), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[5][19] ), .B2(n3144), .Z(n5501) );
  aoim22d1 U4535 ( .A1(n3146), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[5][18] ), .B2(n3144), .Z(n5500) );
  aoim22d1 U4536 ( .A1(n3146), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[5][17] ), .B2(n3143), .Z(n5499) );
  aoim22d1 U4537 ( .A1(n3143), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[5][16] ), .B2(n3143), .Z(n5498) );
  aoim22d1 U4538 ( .A1(n3146), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[5][15] ), .B2(n3143), .Z(n5497) );
  aoim22d1 U4539 ( .A1(n3144), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[5][14] ), .B2(n3143), .Z(n5496) );
  aoim22d1 U4540 ( .A1(n3145), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[5][13] ), .B2(n3143), .Z(n5495) );
  aoim22d1 U4541 ( .A1(n3143), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[5][12] ), .B2(n3143), .Z(n5494) );
  aoim22d1 U4542 ( .A1(n3146), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[5][11] ), .B2(n3145), .Z(n5493) );
  aoim22d1 U4543 ( .A1(n3143), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[5][10] ), .B2(n3145), .Z(n5492) );
  aoim22d1 U4544 ( .A1(n3145), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[5][9] ), .B2(n3145), .Z(n5491) );
  aoim22d1 U4545 ( .A1(n3143), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[5][8] ), .B2(n3145), .Z(n5490) );
  aoim22d1 U4546 ( .A1(n3144), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[5][7] ), .B2(n3145), .Z(n5489) );
  aoim22d1 U4547 ( .A1(n3145), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[5][6] ), .B2(n3145), .Z(n5488) );
  aoim22d1 U4548 ( .A1(n3144), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[5][5] ), .B2(n3146), .Z(n5487) );
  aoim22d1 U4549 ( .A1(n3145), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[5][4] ), .B2(n3146), .Z(n5486) );
  aoim22d1 U4550 ( .A1(n3143), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[5][3] ), .B2(n3146), .Z(n5485) );
  aoim22d1 U4551 ( .A1(n3145), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[5][2] ), .B2(n3146), .Z(n5484) );
  aoim22d1 U4552 ( .A1(n3146), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[5][1] ), .B2(n3146), .Z(n5483) );
  buffd1 U4553 ( .I(n3148), .Z(n3149) );
  buffd1 U4554 ( .I(n3148), .Z(n3152) );
  aoim22d1 U4555 ( .A1(n3149), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[4][0] ), .B2(n3152), .Z(n5482) );
  aoim22d1 U4556 ( .A1(n3152), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[4][31] ), .B2(n3152), .Z(n5481) );
  buffd1 U4557 ( .I(n3148), .Z(n3151) );
  aoim22d1 U4558 ( .A1(n3149), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[4][30] ), .B2(n3151), .Z(n5480) );
  aoim22d1 U4559 ( .A1(n3149), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[4][29] ), .B2(n3151), .Z(n5479) );
  aoim22d1 U4560 ( .A1(n3151), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[4][28] ), .B2(n3151), .Z(n5478) );
  buffd1 U4561 ( .I(n3148), .Z(n3150) );
  aoim22d1 U4562 ( .A1(n3149), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[4][27] ), .B2(n3150), .Z(n5477) );
  aoim22d1 U4563 ( .A1(n3149), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[4][26] ), .B2(n3151), .Z(n5476) );
  aoim22d1 U4564 ( .A1(n3152), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[4][25] ), .B2(n3150), .Z(n5475) );
  aoim22d1 U4565 ( .A1(n3149), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[4][24] ), .B2(n3149), .Z(n5474) );
  aoim22d1 U4566 ( .A1(n3150), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[4][23] ), .B2(n3150), .Z(n5473) );
  aoim22d1 U4567 ( .A1(n3149), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[4][22] ), .B2(n3149), .Z(n5472) );
  aoim22d1 U4568 ( .A1(n3152), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[4][21] ), .B2(n3149), .Z(n5471) );
  aoim22d1 U4569 ( .A1(n3149), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[4][20] ), .B2(n3150), .Z(n5470) );
  aoim22d1 U4570 ( .A1(n3152), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[4][19] ), .B2(n3149), .Z(n5469) );
  aoim22d1 U4571 ( .A1(n3152), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[4][18] ), .B2(n3149), .Z(n5468) );
  aoim22d1 U4572 ( .A1(n3152), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[4][17] ), .B2(n3150), .Z(n5467) );
  aoim22d1 U4573 ( .A1(n3150), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[4][16] ), .B2(n3150), .Z(n5466) );
  aoim22d1 U4574 ( .A1(n3152), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[4][15] ), .B2(n3150), .Z(n5465) );
  aoim22d1 U4575 ( .A1(n3149), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[4][14] ), .B2(n3150), .Z(n5464) );
  aoim22d1 U4576 ( .A1(n3151), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[4][13] ), .B2(n3150), .Z(n5463) );
  aoim22d1 U4577 ( .A1(n3150), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[4][12] ), .B2(n3150), .Z(n5462) );
  aoim22d1 U4578 ( .A1(n3152), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[4][11] ), .B2(n3151), .Z(n5461) );
  aoim22d1 U4579 ( .A1(n3150), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[4][10] ), .B2(n3151), .Z(n5460) );
  aoim22d1 U4580 ( .A1(n3151), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[4][9] ), .B2(n3151), .Z(n5459) );
  aoim22d1 U4581 ( .A1(n3150), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[4][8] ), .B2(n3151), .Z(n5458) );
  aoim22d1 U4582 ( .A1(n3149), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[4][7] ), .B2(n3151), .Z(n5457) );
  aoim22d1 U4583 ( .A1(n3151), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[4][6] ), .B2(n3151), .Z(n5456) );
  aoim22d1 U4584 ( .A1(n3149), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[4][5] ), .B2(n3152), .Z(n5455) );
  aoim22d1 U4585 ( .A1(n3151), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[4][4] ), .B2(n3152), .Z(n5454) );
  aoim22d1 U4586 ( .A1(n3150), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[4][3] ), .B2(n3152), .Z(n5453) );
  aoim22d1 U4587 ( .A1(n3151), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[4][2] ), .B2(n3152), .Z(n5452) );
  aoim22d1 U4588 ( .A1(n3152), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[4][1] ), .B2(n3152), .Z(n5451) );
  nr03d0 U4589 ( .A1(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[2] ), 
        .A2(n3159), .A3(n3165), .ZN(n3154) );
  buffd1 U4590 ( .I(n3154), .Z(n3157) );
  buffd1 U4591 ( .I(n3154), .Z(n3156) );
  aoim22d1 U4592 ( .A1(n3157), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[3][0] ), .B2(n3156), .Z(n5450) );
  aoim22d1 U4593 ( .A1(n3156), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[3][31] ), .B2(n3156), .Z(n5449) );
  buffd1 U4594 ( .I(n3154), .Z(n3155) );
  aoim22d1 U4595 ( .A1(n3157), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[3][30] ), .B2(n3155), .Z(n5448) );
  buffd1 U4596 ( .I(n3155), .Z(n3153) );
  aoim22d1 U4597 ( .A1(n3157), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[3][29] ), .B2(n3153), .Z(n5447) );
  aoim22d1 U4598 ( .A1(n3154), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[3][28] ), .B2(n3155), .Z(n5446) );
  aoim22d1 U4599 ( .A1(n3157), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[3][27] ), .B2(n3153), .Z(n5445) );
  aoim22d1 U4600 ( .A1(n3157), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[3][26] ), .B2(n3155), .Z(n5444) );
  aoim22d1 U4601 ( .A1(n3157), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[3][25] ), .B2(n3153), .Z(n5443) );
  aoim22d1 U4602 ( .A1(n3154), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[3][24] ), .B2(n3157), .Z(n5442) );
  aoim22d1 U4603 ( .A1(n3156), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[3][23] ), .B2(n3153), .Z(n5441) );
  aoim22d1 U4604 ( .A1(n3156), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[3][22] ), .B2(n3157), .Z(n5440) );
  aoim22d1 U4605 ( .A1(n3156), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[3][21] ), .B2(n3157), .Z(n5439) );
  aoim22d1 U4606 ( .A1(n3157), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[3][20] ), .B2(n3153), .Z(n5438) );
  aoim22d1 U4607 ( .A1(n3156), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[3][19] ), .B2(n3157), .Z(n5437) );
  aoim22d1 U4608 ( .A1(n3155), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[3][18] ), .B2(n3157), .Z(n5436) );
  aoim22d1 U4609 ( .A1(n3156), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[3][17] ), .B2(n3153), .Z(n5435) );
  aoim22d1 U4610 ( .A1(n3156), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[3][16] ), .B2(n3153), .Z(n5434) );
  aoim22d1 U4611 ( .A1(n3153), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[3][15] ), .B2(n3153), .Z(n5433) );
  aoim22d1 U4612 ( .A1(n3157), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[3][14] ), .B2(n3153), .Z(n5432) );
  aoim22d1 U4613 ( .A1(n3156), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[3][13] ), .B2(n3153), .Z(n5431) );
  aoim22d1 U4614 ( .A1(n3154), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[3][12] ), .B2(n3153), .Z(n5430) );
  aoim22d1 U4615 ( .A1(n3157), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[3][11] ), .B2(n3157), .Z(n5429) );
  aoim22d1 U4616 ( .A1(n3155), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[3][10] ), .B2(n3156), .Z(n5428) );
  aoim22d1 U4617 ( .A1(n3155), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[3][9] ), .B2(n3155), .Z(n5427) );
  aoim22d1 U4618 ( .A1(n3155), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[3][8] ), .B2(n3157), .Z(n5426) );
  aoim22d1 U4619 ( .A1(n3155), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[3][7] ), .B2(n3156), .Z(n5425) );
  aoim22d1 U4620 ( .A1(n3155), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[3][6] ), .B2(n3155), .Z(n5424) );
  aoim22d1 U4621 ( .A1(n3155), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[3][5] ), .B2(n3156), .Z(n5423) );
  aoim22d1 U4622 ( .A1(n3155), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[3][4] ), .B2(n3156), .Z(n5422) );
  aoim22d1 U4623 ( .A1(n3155), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[3][3] ), .B2(n3156), .Z(n5421) );
  aoim22d1 U4624 ( .A1(n3155), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[3][2] ), .B2(n3156), .Z(n5420) );
  aoim22d1 U4625 ( .A1(n3157), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[3][1] ), .B2(n3156), .Z(n5419) );
  nr03d0 U4626 ( .A1(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[2] ), 
        .A2(n3159), .A3(n3158), .ZN(n3161) );
  buffd1 U4627 ( .I(n3161), .Z(n3164) );
  buffd1 U4628 ( .I(n3161), .Z(n3163) );
  aoim22d1 U4629 ( .A1(n3164), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[2][0] ), .B2(n3163), .Z(n5418) );
  aoim22d1 U4630 ( .A1(n3163), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[2][31] ), .B2(n3163), .Z(n5417) );
  buffd1 U4631 ( .I(n3161), .Z(n3162) );
  aoim22d1 U4632 ( .A1(n3164), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[2][30] ), .B2(n3162), .Z(n5416) );
  buffd1 U4633 ( .I(n3162), .Z(n3160) );
  aoim22d1 U4634 ( .A1(n3164), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[2][29] ), .B2(n3160), .Z(n5415) );
  aoim22d1 U4635 ( .A1(n3161), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[2][28] ), .B2(n3162), .Z(n5414) );
  aoim22d1 U4636 ( .A1(n3164), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[2][27] ), .B2(n3160), .Z(n5413) );
  aoim22d1 U4637 ( .A1(n3164), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[2][26] ), .B2(n3162), .Z(n5412) );
  aoim22d1 U4638 ( .A1(n3164), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[2][25] ), .B2(n3160), .Z(n5411) );
  aoim22d1 U4639 ( .A1(n3161), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[2][24] ), .B2(n3164), .Z(n5410) );
  aoim22d1 U4640 ( .A1(n3163), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[2][23] ), .B2(n3160), .Z(n5409) );
  aoim22d1 U4641 ( .A1(n3163), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[2][22] ), .B2(n3164), .Z(n5408) );
  aoim22d1 U4642 ( .A1(n3163), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[2][21] ), .B2(n3164), .Z(n5407) );
  aoim22d1 U4643 ( .A1(n3164), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[2][20] ), .B2(n3160), .Z(n5406) );
  aoim22d1 U4644 ( .A1(n3163), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[2][19] ), .B2(n3164), .Z(n5405) );
  aoim22d1 U4645 ( .A1(n3162), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[2][18] ), .B2(n3164), .Z(n5404) );
  aoim22d1 U4646 ( .A1(n3163), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[2][17] ), .B2(n3160), .Z(n5403) );
  aoim22d1 U4647 ( .A1(n3163), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[2][16] ), .B2(n3160), .Z(n5402) );
  aoim22d1 U4648 ( .A1(n3160), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[2][15] ), .B2(n3160), .Z(n5401) );
  aoim22d1 U4649 ( .A1(n3164), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[2][14] ), .B2(n3160), .Z(n5400) );
  aoim22d1 U4650 ( .A1(n3163), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[2][13] ), .B2(n3160), .Z(n5399) );
  aoim22d1 U4651 ( .A1(n3161), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[2][12] ), .B2(n3160), .Z(n5398) );
  aoim22d1 U4652 ( .A1(n3164), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[2][11] ), .B2(n3164), .Z(n5397) );
  aoim22d1 U4653 ( .A1(n3162), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[2][10] ), .B2(n3163), .Z(n5396) );
  aoim22d1 U4654 ( .A1(n3162), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[2][9] ), .B2(n3162), .Z(n5395) );
  aoim22d1 U4655 ( .A1(n3162), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[2][8] ), .B2(n3164), .Z(n5394) );
  aoim22d1 U4656 ( .A1(n3162), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[2][7] ), .B2(n3163), .Z(n5393) );
  aoim22d1 U4657 ( .A1(n3162), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[2][6] ), .B2(n3162), .Z(n5392) );
  aoim22d1 U4658 ( .A1(n3162), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[2][5] ), .B2(n3163), .Z(n5391) );
  aoim22d1 U4659 ( .A1(n3162), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[2][4] ), .B2(n3163), .Z(n5390) );
  aoim22d1 U4660 ( .A1(n3162), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[2][3] ), .B2(n3163), .Z(n5389) );
  aoim22d1 U4661 ( .A1(n3162), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[2][2] ), .B2(n3163), .Z(n5388) );
  aoim22d1 U4662 ( .A1(n3164), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[2][1] ), .B2(n3163), .Z(n5387) );
  nr03d0 U4663 ( .A1(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[1] ), 
        .A2(
        \IBusCachedPlugin_cache/lineLoader_write_data_0_payload_address[2] ), 
        .A3(n3165), .ZN(n3168) );
  buffd1 U4664 ( .I(n3168), .Z(n3171) );
  buffd1 U4665 ( .I(n3168), .Z(n3170) );
  aoim22d1 U4666 ( .A1(n3171), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[1][0] ), .B2(n3170), .Z(n5386) );
  aoim22d1 U4667 ( .A1(n3170), .A2(n3166), .B1(
        \IBusCachedPlugin_cache/banks_0[1][31] ), .B2(n3170), .Z(n5385) );
  buffd1 U4668 ( .I(n3168), .Z(n3169) );
  aoim22d1 U4669 ( .A1(n3171), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[1][30] ), .B2(n3169), .Z(n5384) );
  buffd1 U4670 ( .I(n3169), .Z(n3167) );
  aoim22d1 U4671 ( .A1(n3171), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[1][29] ), .B2(n3167), .Z(n5383) );
  aoim22d1 U4672 ( .A1(n3168), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[1][28] ), .B2(n3169), .Z(n5382) );
  aoim22d1 U4673 ( .A1(n3171), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[1][27] ), .B2(n3167), .Z(n5381) );
  aoim22d1 U4674 ( .A1(n3171), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[1][26] ), .B2(n3169), .Z(n5380) );
  aoim22d1 U4675 ( .A1(n3171), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[1][25] ), .B2(n3167), .Z(n5379) );
  aoim22d1 U4676 ( .A1(n3168), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[1][24] ), .B2(n3171), .Z(n5378) );
  aoim22d1 U4677 ( .A1(n3170), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[1][23] ), .B2(n3167), .Z(n5377) );
  aoim22d1 U4678 ( .A1(n3170), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[1][22] ), .B2(n3171), .Z(n5376) );
  aoim22d1 U4679 ( .A1(n3170), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[1][21] ), .B2(n3171), .Z(n5375) );
  aoim22d1 U4680 ( .A1(n3171), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[1][20] ), .B2(n3167), .Z(n5374) );
  aoim22d1 U4681 ( .A1(n3170), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[1][19] ), .B2(n3171), .Z(n5373) );
  aoim22d1 U4682 ( .A1(n3169), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[1][18] ), .B2(n3171), .Z(n5372) );
  aoim22d1 U4683 ( .A1(n3170), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[1][17] ), .B2(n3167), .Z(n5371) );
  aoim22d1 U4684 ( .A1(n3170), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[1][16] ), .B2(n3167), .Z(n5370) );
  aoim22d1 U4685 ( .A1(n3167), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[1][15] ), .B2(n3167), .Z(n5369) );
  aoim22d1 U4686 ( .A1(n3171), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[1][14] ), .B2(n3167), .Z(n5368) );
  aoim22d1 U4687 ( .A1(n3170), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[1][13] ), .B2(n3167), .Z(n5367) );
  aoim22d1 U4688 ( .A1(n3168), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[1][12] ), .B2(n3167), .Z(n5366) );
  aoim22d1 U4689 ( .A1(n3171), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[1][11] ), .B2(n3171), .Z(n5365) );
  aoim22d1 U4690 ( .A1(n3169), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[1][10] ), .B2(n3170), .Z(n5364) );
  aoim22d1 U4691 ( .A1(n3169), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[1][9] ), .B2(n3169), .Z(n5363) );
  aoim22d1 U4692 ( .A1(n3169), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[1][8] ), .B2(n3171), .Z(n5362) );
  aoim22d1 U4693 ( .A1(n3169), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[1][7] ), .B2(n3170), .Z(n5361) );
  aoim22d1 U4694 ( .A1(n3169), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[1][6] ), .B2(n3169), .Z(n5360) );
  aoim22d1 U4695 ( .A1(n3169), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[1][5] ), .B2(n3170), .Z(n5359) );
  aoim22d1 U4696 ( .A1(n3169), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[1][4] ), .B2(n3170), .Z(n5358) );
  aoim22d1 U4697 ( .A1(n3169), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[1][3] ), .B2(n3170), .Z(n5357) );
  aoim22d1 U4698 ( .A1(n3169), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[1][2] ), .B2(n3170), .Z(n5356) );
  aoim22d1 U4699 ( .A1(n3171), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[1][1] ), .B2(n3170), .Z(n5355) );
  aoim22d1 U4700 ( .A1(n3207), .A2(n3172), .B1(
        \IBusCachedPlugin_cache/banks_0[0][0] ), .B2(n3207), .Z(n5354) );
  buffd1 U4701 ( .I(n3191), .Z(n3205) );
  aoim22d1 U4702 ( .A1(n3197), .A2(n3173), .B1(
        \IBusCachedPlugin_cache/banks_0[0][30] ), .B2(n3205), .Z(n5353) );
  buffd1 U4703 ( .I(n3205), .Z(n3192) );
  aoim22d1 U4704 ( .A1(n3197), .A2(n3174), .B1(
        \IBusCachedPlugin_cache/banks_0[0][29] ), .B2(n3192), .Z(n5352) );
  aoim22d1 U4705 ( .A1(n3191), .A2(n3175), .B1(
        \IBusCachedPlugin_cache/banks_0[0][28] ), .B2(n3205), .Z(n5351) );
  aoim22d1 U4706 ( .A1(n3197), .A2(n3176), .B1(
        \IBusCachedPlugin_cache/banks_0[0][27] ), .B2(n3192), .Z(n5350) );
  aoim22d1 U4707 ( .A1(n3197), .A2(n3177), .B1(
        \IBusCachedPlugin_cache/banks_0[0][26] ), .B2(n3205), .Z(n5349) );
  aoim22d1 U4708 ( .A1(n3197), .A2(n3178), .B1(
        \IBusCachedPlugin_cache/banks_0[0][25] ), .B2(n3192), .Z(n5348) );
  aoim22d1 U4709 ( .A1(n3191), .A2(n3179), .B1(
        \IBusCachedPlugin_cache/banks_0[0][24] ), .B2(n3197), .Z(n5347) );
  aoim22d1 U4710 ( .A1(n3207), .A2(n3180), .B1(
        \IBusCachedPlugin_cache/banks_0[0][23] ), .B2(n3192), .Z(n5346) );
  aoim22d1 U4711 ( .A1(n3207), .A2(n3181), .B1(
        \IBusCachedPlugin_cache/banks_0[0][22] ), .B2(n3197), .Z(n5345) );
  aoim22d1 U4712 ( .A1(n3197), .A2(n3182), .B1(
        \IBusCachedPlugin_cache/banks_0[0][21] ), .B2(n3197), .Z(n5344) );
  aoim22d1 U4713 ( .A1(n3207), .A2(n3183), .B1(
        \IBusCachedPlugin_cache/banks_0[0][20] ), .B2(n3192), .Z(n5343) );
  aoim22d1 U4714 ( .A1(n3205), .A2(n3184), .B1(
        \IBusCachedPlugin_cache/banks_0[0][19] ), .B2(n3197), .Z(n5342) );
  aoim22d1 U4715 ( .A1(n3197), .A2(n3185), .B1(
        \IBusCachedPlugin_cache/banks_0[0][18] ), .B2(n3197), .Z(n5341) );
  aoim22d1 U4716 ( .A1(n3207), .A2(n3186), .B1(
        \IBusCachedPlugin_cache/banks_0[0][17] ), .B2(n3192), .Z(n5340) );
  aoim22d1 U4717 ( .A1(n3192), .A2(n3187), .B1(
        \IBusCachedPlugin_cache/banks_0[0][16] ), .B2(n3192), .Z(n5339) );
  aoim22d1 U4718 ( .A1(n3197), .A2(n3188), .B1(
        \IBusCachedPlugin_cache/banks_0[0][15] ), .B2(n3192), .Z(n5338) );
  aoim22d1 U4719 ( .A1(n3207), .A2(n3189), .B1(
        \IBusCachedPlugin_cache/banks_0[0][14] ), .B2(n3192), .Z(n5337) );
  aoim22d1 U4720 ( .A1(n3191), .A2(n3190), .B1(
        \IBusCachedPlugin_cache/banks_0[0][13] ), .B2(n3192), .Z(n5336) );
  aoim22d1 U4721 ( .A1(n3197), .A2(n3193), .B1(
        \IBusCachedPlugin_cache/banks_0[0][12] ), .B2(n3192), .Z(n5335) );
  aoim22d1 U4722 ( .A1(n3207), .A2(n3194), .B1(
        \IBusCachedPlugin_cache/banks_0[0][11] ), .B2(n3197), .Z(n5334) );
  aoim22d1 U4723 ( .A1(n3205), .A2(n3195), .B1(
        \IBusCachedPlugin_cache/banks_0[0][10] ), .B2(n3207), .Z(n5333) );
  aoim22d1 U4724 ( .A1(n3205), .A2(n3196), .B1(
        \IBusCachedPlugin_cache/banks_0[0][9] ), .B2(n3205), .Z(n5332) );
  aoim22d1 U4725 ( .A1(n3205), .A2(n3198), .B1(
        \IBusCachedPlugin_cache/banks_0[0][8] ), .B2(n3197), .Z(n5331) );
  aoim22d1 U4726 ( .A1(n3205), .A2(n3199), .B1(
        \IBusCachedPlugin_cache/banks_0[0][7] ), .B2(n3207), .Z(n5330) );
  aoim22d1 U4727 ( .A1(n3205), .A2(n3200), .B1(
        \IBusCachedPlugin_cache/banks_0[0][6] ), .B2(n3205), .Z(n5329) );
  aoim22d1 U4728 ( .A1(n3205), .A2(n3201), .B1(
        \IBusCachedPlugin_cache/banks_0[0][5] ), .B2(n3207), .Z(n5328) );
  aoim22d1 U4729 ( .A1(n3205), .A2(n3202), .B1(
        \IBusCachedPlugin_cache/banks_0[0][4] ), .B2(n3207), .Z(n5327) );
  aoim22d1 U4730 ( .A1(n3205), .A2(n3203), .B1(
        \IBusCachedPlugin_cache/banks_0[0][3] ), .B2(n3207), .Z(n5326) );
  aoim22d1 U4731 ( .A1(n3205), .A2(n3204), .B1(
        \IBusCachedPlugin_cache/banks_0[0][2] ), .B2(n3207), .Z(n5325) );
  aoim22d1 U4732 ( .A1(n3207), .A2(n3206), .B1(
        \IBusCachedPlugin_cache/banks_0[0][1] ), .B2(n3207), .Z(n5324) );
  inv0d0 U4733 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[31]), .ZN(
        n3824) );
  inv0d0 U4734 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[31]), .ZN(
        n3208) );
  aoi22d1 U4735 ( .A1(n6893), .A2(n3824), .B1(n3208), .B2(n6908), .ZN(n5318)
         );
  aoi22d1 U4736 ( .A1(n3209), .A2(n3208), .B1(n6416), .B2(n3232), .ZN(n5317)
         );
  inv0d0 U4737 ( .I(writeBack_PC[31]), .ZN(n3663) );
  inv0d0 U4738 ( .I(memory_PC[31]), .ZN(n6417) );
  aoi22d1 U4739 ( .A1(CsrPlugin_exceptionPendings_3), .A2(n3663), .B1(n6417), 
        .B2(n3245), .ZN(n5316) );
  inv0d0 U4740 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[30]), .ZN(
        n3822) );
  inv0d0 U4741 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[30]), .ZN(
        n3210) );
  aoi22d1 U4742 ( .A1(n6893), .A2(n3822), .B1(n3210), .B2(n6908), .ZN(n5315)
         );
  aoi22d1 U4743 ( .A1(n3249), .A2(n3210), .B1(n6418), .B2(n3243), .ZN(n5314)
         );
  inv0d0 U4744 ( .I(writeBack_PC[30]), .ZN(n3657) );
  inv0d0 U4745 ( .I(memory_PC[30]), .ZN(n6419) );
  aoi22d1 U4746 ( .A1(CsrPlugin_exceptionPendings_3), .A2(n3657), .B1(n6419), 
        .B2(n3245), .ZN(n5313) );
  inv0d0 U4747 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[29]), .ZN(
        n6808) );
  inv0d0 U4748 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[29]), .ZN(
        n3211) );
  aoi22d1 U4749 ( .A1(n6893), .A2(n6808), .B1(n3211), .B2(n6936), .ZN(n5312)
         );
  aoi22d1 U4750 ( .A1(n3249), .A2(n3211), .B1(n6809), .B2(n3243), .ZN(n5311)
         );
  inv0d0 U4751 ( .I(writeBack_PC[29]), .ZN(n3653) );
  inv0d0 U4752 ( .I(memory_PC[29]), .ZN(n6810) );
  aoi22d1 U4753 ( .A1(CsrPlugin_exceptionPendings_3), .A2(n3653), .B1(n6810), 
        .B2(n3245), .ZN(n5310) );
  inv0d0 U4754 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[28]), .ZN(
        n6813) );
  inv0d0 U4755 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[28]), .ZN(
        n3212) );
  aoi22d1 U4756 ( .A1(n6893), .A2(n6813), .B1(n3212), .B2(n6936), .ZN(n5309)
         );
  aoi22d1 U4757 ( .A1(n3249), .A2(n3212), .B1(n6814), .B2(n3247), .ZN(n5308)
         );
  inv0d0 U4758 ( .I(writeBack_PC[28]), .ZN(n3650) );
  inv0d0 U4759 ( .I(memory_PC[28]), .ZN(n6815) );
  aoi22d1 U4760 ( .A1(n3230), .A2(n3650), .B1(n6815), .B2(n3245), .ZN(n5307)
         );
  inv0d0 U4761 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[27]), .ZN(
        n6818) );
  inv0d0 U4762 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[27]), .ZN(
        n3213) );
  aoi22d1 U4763 ( .A1(n6893), .A2(n6818), .B1(n3213), .B2(n6936), .ZN(n5306)
         );
  aoi22d1 U4764 ( .A1(n3249), .A2(n3213), .B1(n6819), .B2(n3232), .ZN(n5305)
         );
  inv0d0 U4765 ( .I(writeBack_PC[27]), .ZN(n3647) );
  inv0d0 U4766 ( .I(memory_PC[27]), .ZN(n6820) );
  aoi22d1 U4767 ( .A1(n3230), .A2(n3647), .B1(n6820), .B2(n3245), .ZN(n5304)
         );
  inv0d0 U4768 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[26]), .ZN(
        n6823) );
  inv0d0 U4769 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[26]), .ZN(
        n3214) );
  aoi22d1 U4770 ( .A1(n6893), .A2(n6823), .B1(n3214), .B2(n6862), .ZN(n5303)
         );
  aoi22d1 U4771 ( .A1(n3249), .A2(n3214), .B1(n6824), .B2(n3247), .ZN(n5302)
         );
  inv0d0 U4772 ( .I(writeBack_PC[26]), .ZN(n3644) );
  inv0d0 U4773 ( .I(memory_PC[26]), .ZN(n6825) );
  aoi22d1 U4774 ( .A1(n3230), .A2(n3644), .B1(n6825), .B2(n3245), .ZN(n5301)
         );
  inv0d0 U4775 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[25]), .ZN(
        n6828) );
  inv0d0 U4776 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[25]), .ZN(
        n3215) );
  aoi22d1 U4777 ( .A1(n6893), .A2(n6828), .B1(n3215), .B2(n6862), .ZN(n5300)
         );
  aoi22d1 U4778 ( .A1(n3249), .A2(n3215), .B1(n6829), .B2(n3247), .ZN(n5299)
         );
  inv0d0 U4779 ( .I(writeBack_PC[25]), .ZN(n3640) );
  inv0d0 U4780 ( .I(memory_PC[25]), .ZN(n6830) );
  aoi22d1 U4781 ( .A1(n3230), .A2(n3640), .B1(n6830), .B2(n3250), .ZN(n5298)
         );
  inv0d0 U4782 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[24]), .ZN(
        n6833) );
  inv0d0 U4783 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[24]), .ZN(
        n3216) );
  buffd1 U4784 ( .I(n6862), .Z(n6999) );
  aoi22d1 U4785 ( .A1(n6893), .A2(n6833), .B1(n3216), .B2(n6999), .ZN(n5297)
         );
  aoi22d1 U4786 ( .A1(n3249), .A2(n3216), .B1(n6834), .B2(n3243), .ZN(n5296)
         );
  inv0d0 U4787 ( .I(writeBack_PC[24]), .ZN(n3639) );
  inv0d0 U4788 ( .I(memory_PC[24]), .ZN(n6835) );
  aoi22d1 U4789 ( .A1(n3230), .A2(n3639), .B1(n6835), .B2(n3245), .ZN(n5295)
         );
  inv0d0 U4790 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[23]), .ZN(
        n6838) );
  inv0d0 U4791 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[23]), .ZN(
        n3217) );
  aoi22d1 U4792 ( .A1(n6893), .A2(n6838), .B1(n3217), .B2(n6999), .ZN(n5294)
         );
  aoi22d1 U4793 ( .A1(n3249), .A2(n3217), .B1(n6839), .B2(n3232), .ZN(n5293)
         );
  inv0d0 U4794 ( .I(writeBack_PC[23]), .ZN(n3634) );
  inv0d0 U4795 ( .I(memory_PC[23]), .ZN(n6840) );
  aoi22d1 U4796 ( .A1(n3230), .A2(n3634), .B1(n6840), .B2(n3250), .ZN(n5292)
         );
  inv0d0 U4797 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[22]), .ZN(
        n6843) );
  inv0d0 U4798 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[22]), .ZN(
        n3218) );
  aoi22d1 U4799 ( .A1(n6893), .A2(n6843), .B1(n3218), .B2(n6862), .ZN(n5291)
         );
  aoi22d1 U4800 ( .A1(n3249), .A2(n3218), .B1(n6844), .B2(n3232), .ZN(n5290)
         );
  inv0d0 U4801 ( .I(writeBack_PC[22]), .ZN(n3633) );
  inv0d0 U4802 ( .I(memory_PC[22]), .ZN(n6845) );
  aoi22d1 U4803 ( .A1(n3230), .A2(n3633), .B1(n6845), .B2(n3250), .ZN(n5289)
         );
  inv0d0 U4804 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[21]), .ZN(
        n6848) );
  inv0d0 U4805 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[21]), .ZN(
        n3219) );
  aoi22d1 U4806 ( .A1(n6893), .A2(n6848), .B1(n3219), .B2(n6936), .ZN(n5288)
         );
  aoi22d1 U4807 ( .A1(n3249), .A2(n3219), .B1(n6849), .B2(n3232), .ZN(n5287)
         );
  inv0d0 U4808 ( .I(writeBack_PC[21]), .ZN(n3628) );
  inv0d0 U4809 ( .I(memory_PC[21]), .ZN(n6850) );
  aoi22d1 U4810 ( .A1(n3230), .A2(n3628), .B1(n6850), .B2(n3245), .ZN(n5286)
         );
  inv0d0 U4811 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[20]), .ZN(
        n6853) );
  inv0d0 U4812 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[20]), .ZN(
        n3220) );
  aoi22d1 U4813 ( .A1(n6893), .A2(n6853), .B1(n3220), .B2(n6862), .ZN(n5285)
         );
  aoi22d1 U4814 ( .A1(n3559), .A2(n3220), .B1(n6854), .B2(n3232), .ZN(n5284)
         );
  inv0d0 U4815 ( .I(writeBack_PC[20]), .ZN(n3625) );
  inv0d0 U4816 ( .I(memory_PC[20]), .ZN(n6855) );
  aoi22d1 U4817 ( .A1(n3230), .A2(n3625), .B1(n6855), .B2(n3245), .ZN(n5283)
         );
  inv0d0 U4818 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[19]), .ZN(
        n6858) );
  inv0d0 U4819 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[19]), .ZN(
        n3221) );
  aoi22d1 U4820 ( .A1(n6893), .A2(n6858), .B1(n3221), .B2(n6862), .ZN(n5282)
         );
  aoi22d1 U4821 ( .A1(n3559), .A2(n3221), .B1(n6859), .B2(n3232), .ZN(n5281)
         );
  inv0d0 U4822 ( .I(writeBack_PC[19]), .ZN(n3622) );
  inv0d0 U4823 ( .I(memory_PC[19]), .ZN(n6860) );
  aoi22d1 U4824 ( .A1(n3230), .A2(n3622), .B1(n6860), .B2(n3250), .ZN(n5280)
         );
  inv0d0 U4825 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[18]), .ZN(
        n6864) );
  inv0d0 U4826 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[18]), .ZN(
        n3222) );
  aoi22d1 U4827 ( .A1(n6893), .A2(n6864), .B1(n3222), .B2(n6936), .ZN(n5279)
         );
  aoi22d1 U4828 ( .A1(n3559), .A2(n3222), .B1(n6865), .B2(n3232), .ZN(n5278)
         );
  inv0d0 U4829 ( .I(writeBack_PC[18]), .ZN(n3619) );
  inv0d0 U4830 ( .I(memory_PC[18]), .ZN(n6866) );
  aoi22d1 U4831 ( .A1(n3230), .A2(n3619), .B1(n6866), .B2(n3250), .ZN(n5277)
         );
  inv0d0 U4832 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[17]), .ZN(
        n6869) );
  inv0d0 U4833 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[17]), .ZN(
        n3223) );
  aoi22d1 U4834 ( .A1(n6893), .A2(n6869), .B1(n3223), .B2(n6999), .ZN(n5276)
         );
  aoi22d1 U4835 ( .A1(n3559), .A2(n3223), .B1(n6870), .B2(n3232), .ZN(n5275)
         );
  inv0d0 U4836 ( .I(writeBack_PC[17]), .ZN(n3616) );
  inv0d0 U4837 ( .I(memory_PC[17]), .ZN(n6871) );
  aoi22d1 U4838 ( .A1(n3230), .A2(n3616), .B1(n6871), .B2(n3250), .ZN(n5274)
         );
  inv0d0 U4839 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[16]), .ZN(
        n6874) );
  inv0d0 U4840 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[16]), .ZN(
        n3224) );
  aoi22d1 U4841 ( .A1(n6893), .A2(n6874), .B1(n3224), .B2(n6999), .ZN(n5273)
         );
  aoi22d1 U4842 ( .A1(n3559), .A2(n3224), .B1(n6875), .B2(n3247), .ZN(n5272)
         );
  inv0d0 U4843 ( .I(writeBack_PC[16]), .ZN(n3613) );
  inv0d0 U4844 ( .I(memory_PC[16]), .ZN(n6876) );
  aoi22d1 U4845 ( .A1(n3230), .A2(n3613), .B1(n6876), .B2(n3250), .ZN(n5271)
         );
  inv0d2 U4846 ( .I(n6936), .ZN(n7090) );
  inv0d0 U4847 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[15]), .ZN(
        n6881) );
  inv0d0 U4848 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[15]), .ZN(
        n3225) );
  aoi22d1 U4849 ( .A1(n7090), .A2(n6881), .B1(n3225), .B2(n6862), .ZN(n5270)
         );
  aoi22d1 U4850 ( .A1(n3559), .A2(n3225), .B1(n6882), .B2(n3243), .ZN(n5269)
         );
  inv0d0 U4851 ( .I(writeBack_PC[15]), .ZN(n3610) );
  inv0d0 U4852 ( .I(memory_PC[15]), .ZN(n6883) );
  aoi22d1 U4853 ( .A1(n3230), .A2(n3610), .B1(n6883), .B2(n3250), .ZN(n5268)
         );
  inv0d0 U4854 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[14]), .ZN(
        n6886) );
  inv0d0 U4855 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[14]), .ZN(
        n3226) );
  aoi22d1 U4856 ( .A1(n7090), .A2(n6886), .B1(n3226), .B2(n6999), .ZN(n5267)
         );
  aoi22d1 U4857 ( .A1(n3559), .A2(n3226), .B1(n6887), .B2(n3243), .ZN(n5266)
         );
  inv0d0 U4858 ( .I(writeBack_PC[14]), .ZN(n3607) );
  inv0d0 U4859 ( .I(memory_PC[14]), .ZN(n6888) );
  aoi22d1 U4860 ( .A1(n3230), .A2(n3607), .B1(n6888), .B2(n3250), .ZN(n5265)
         );
  inv0d0 U4861 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[13]), .ZN(
        n6892) );
  inv0d0 U4862 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[13]), .ZN(
        n3227) );
  aoi22d1 U4863 ( .A1(n6893), .A2(n6892), .B1(n3227), .B2(n6999), .ZN(n5264)
         );
  aoi22d1 U4864 ( .A1(n3559), .A2(n3227), .B1(n6894), .B2(n3247), .ZN(n5263)
         );
  inv0d0 U4865 ( .I(writeBack_PC[13]), .ZN(n3604) );
  inv0d0 U4866 ( .I(memory_PC[13]), .ZN(n6895) );
  aoi22d1 U4867 ( .A1(n3230), .A2(n3604), .B1(n6895), .B2(n3250), .ZN(n5262)
         );
  inv0d0 U4868 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[12]), .ZN(
        n3820) );
  inv0d0 U4869 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[12]), .ZN(
        n3228) );
  aoi22d1 U4870 ( .A1(n7090), .A2(n3820), .B1(n3228), .B2(n6999), .ZN(n5261)
         );
  aoi22d1 U4871 ( .A1(n3559), .A2(n3228), .B1(n7118), .B2(n3243), .ZN(n5260)
         );
  inv0d0 U4872 ( .I(writeBack_PC[12]), .ZN(n3601) );
  inv0d0 U4873 ( .I(memory_PC[12]), .ZN(n7119) );
  aoi22d1 U4874 ( .A1(n3230), .A2(n3601), .B1(n7119), .B2(n3250), .ZN(n5259)
         );
  inv0d0 U4875 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[11]), .ZN(
        n6899) );
  inv0d0 U4876 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[11]), .ZN(
        n3229) );
  aoi22d1 U4877 ( .A1(n7090), .A2(n6899), .B1(n3229), .B2(n6999), .ZN(n5258)
         );
  aoi22d1 U4878 ( .A1(n3559), .A2(n3229), .B1(n6900), .B2(n3247), .ZN(n5257)
         );
  inv0d0 U4879 ( .I(writeBack_PC[11]), .ZN(n3598) );
  inv0d0 U4880 ( .I(memory_PC[11]), .ZN(n6901) );
  aoi22d1 U4881 ( .A1(n3230), .A2(n3598), .B1(n6901), .B2(n3250), .ZN(n5256)
         );
  inv0d0 U4882 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[10]), .ZN(
        n6904) );
  inv0d0 U4883 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[10]), .ZN(
        n3231) );
  aoi22d1 U4884 ( .A1(n7090), .A2(n6904), .B1(n3231), .B2(n6999), .ZN(n5255)
         );
  aoi22d1 U4885 ( .A1(n3559), .A2(n3231), .B1(n6905), .B2(n3232), .ZN(n5254)
         );
  inv0d0 U4886 ( .I(writeBack_PC[10]), .ZN(n3595) );
  inv0d0 U4887 ( .I(memory_PC[10]), .ZN(n6906) );
  aoi22d1 U4888 ( .A1(CsrPlugin_exceptionPendings_3), .A2(n3595), .B1(n6906), 
        .B2(n3250), .ZN(n5253) );
  inv0d0 U4889 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[9]), .ZN(
        n6910) );
  inv0d0 U4890 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[9]), .ZN(
        n3233) );
  aoi22d1 U4891 ( .A1(n7090), .A2(n6910), .B1(n3233), .B2(n6999), .ZN(n5252)
         );
  aoi22d1 U4892 ( .A1(n3559), .A2(n3233), .B1(n6911), .B2(n3232), .ZN(n5251)
         );
  inv0d0 U4893 ( .I(writeBack_PC[9]), .ZN(n3592) );
  inv0d0 U4894 ( .I(memory_PC[9]), .ZN(n6912) );
  aoi22d1 U4895 ( .A1(CsrPlugin_exceptionPendings_3), .A2(n3592), .B1(n6912), 
        .B2(n3250), .ZN(n5250) );
  inv0d0 U4896 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[8]), .ZN(
        n6915) );
  inv0d0 U4897 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[8]), .ZN(
        n3234) );
  aoi22d1 U4898 ( .A1(n7090), .A2(n6915), .B1(n3234), .B2(n6999), .ZN(n5249)
         );
  aoi22d1 U4899 ( .A1(n3559), .A2(n3234), .B1(n6916), .B2(n3235), .ZN(n5248)
         );
  inv0d0 U4900 ( .I(writeBack_PC[8]), .ZN(n3589) );
  inv0d0 U4901 ( .I(memory_PC[8]), .ZN(n6917) );
  aoi22d1 U4902 ( .A1(CsrPlugin_exceptionPendings_3), .A2(n3589), .B1(n6917), 
        .B2(n3245), .ZN(n5247) );
  inv0d0 U4903 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[7]), .ZN(
        n6925) );
  inv0d0 U4904 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[7]), .ZN(
        n3236) );
  aoi22d1 U4905 ( .A1(n7090), .A2(n6925), .B1(n3236), .B2(n6999), .ZN(n5246)
         );
  aoi22d1 U4906 ( .A1(n3559), .A2(n3236), .B1(n6927), .B2(n3235), .ZN(n5245)
         );
  inv0d0 U4907 ( .I(writeBack_PC[7]), .ZN(n3586) );
  inv0d0 U4908 ( .I(memory_PC[7]), .ZN(n6928) );
  aoi22d1 U4909 ( .A1(CsrPlugin_exceptionPendings_3), .A2(n3586), .B1(n6928), 
        .B2(n3245), .ZN(n5244) );
  inv0d0 U4910 ( .I(IBusCachedPlugin_iBusRsp_stages_1_input_payload[6]), .ZN(
        n6938) );
  inv0d0 U4911 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[6]), .ZN(
        n3237) );
  aoi22d1 U4912 ( .A1(n7090), .A2(n6938), .B1(n3237), .B2(n6999), .ZN(n5243)
         );
  aoi22d1 U4913 ( .A1(n3249), .A2(n3237), .B1(n6940), .B2(n3243), .ZN(n5242)
         );
  inv0d0 U4914 ( .I(writeBack_PC[6]), .ZN(n3583) );
  inv0d0 U4915 ( .I(memory_PC[6]), .ZN(n6941) );
  aoi22d1 U4916 ( .A1(CsrPlugin_exceptionPendings_3), .A2(n3583), .B1(n6941), 
        .B2(n3245), .ZN(n5241) );
  inv0d1 U4917 ( .I(n6936), .ZN(n7085) );
  inv0d0 U4918 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[5]), .ZN(
        n3239) );
  aoi22d1 U4919 ( .A1(n7085), .A2(n7001), .B1(n3239), .B2(n6999), .ZN(n5240)
         );
  aoi22d1 U4920 ( .A1(n3249), .A2(n3239), .B1(n7002), .B2(n3238), .ZN(n5239)
         );
  inv0d0 U4921 ( .I(writeBack_PC[5]), .ZN(n3580) );
  inv0d0 U4922 ( .I(memory_PC[5]), .ZN(n7003) );
  aoi22d1 U4923 ( .A1(CsrPlugin_exceptionPendings_3), .A2(n3580), .B1(n7003), 
        .B2(n3245), .ZN(n5238) );
  inv0d0 U4924 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[4]), .ZN(
        n3241) );
  aoi22d1 U4925 ( .A1(n7090), .A2(n3240), .B1(n3241), .B2(n6999), .ZN(n5237)
         );
  aoi22d1 U4926 ( .A1(n3559), .A2(n3241), .B1(n7114), .B2(n3243), .ZN(n5236)
         );
  inv0d0 U4927 ( .I(writeBack_PC[4]), .ZN(n3577) );
  inv0d0 U4928 ( .I(memory_PC[4]), .ZN(n7115) );
  aoi22d1 U4929 ( .A1(CsrPlugin_exceptionPendings_3), .A2(n3577), .B1(n7115), 
        .B2(n3245), .ZN(n5235) );
  inv0d1 U4930 ( .I(n6908), .ZN(n6939) );
  inv0d0 U4931 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[3]), .ZN(
        n3244) );
  aoi22d1 U4932 ( .A1(n6939), .A2(n3242), .B1(n3244), .B2(n6999), .ZN(n5234)
         );
  aoi22d1 U4933 ( .A1(n3249), .A2(n3244), .B1(n6420), .B2(n3243), .ZN(n5233)
         );
  inv0d0 U4934 ( .I(writeBack_PC[3]), .ZN(n3574) );
  inv0d0 U4935 ( .I(memory_PC[3]), .ZN(n6421) );
  aoi22d1 U4936 ( .A1(CsrPlugin_exceptionPendings_3), .A2(n3574), .B1(n6421), 
        .B2(n3245), .ZN(n5232) );
  inv0d0 U4937 ( .I(
        IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload[2]), .ZN(
        n3248) );
  aoi22d1 U4938 ( .A1(n6939), .A2(n3246), .B1(n3248), .B2(n6862), .ZN(n5231)
         );
  aoi22d1 U4939 ( .A1(n3249), .A2(n3248), .B1(n6299), .B2(n3247), .ZN(n5230)
         );
  inv0d0 U4940 ( .I(writeBack_PC[2]), .ZN(n3571) );
  inv0d0 U4941 ( .I(memory_PC[2]), .ZN(n3825) );
  aoi22d1 U4942 ( .A1(CsrPlugin_exceptionPendings_3), .A2(n3571), .B1(n3825), 
        .B2(n3250), .ZN(n5229) );
  nr02d0 U4943 ( .A1(n3316), .A2(n3287), .ZN(n3309) );
  nd03d0 U4944 ( .A1(_zz_lastStageRegFileWrite_payload_address[9]), .A2(
        _zz_lastStageRegFileWrite_payload_address[8]), .A3(n3309), .ZN(n3434)
         );
  nd04d0 U4945 ( .A1(_zz_lastStageRegFileWrite_payload_address[10]), .A2(
        _zz_lastStageRegFileWrite_payload_address[11]), .A3(n3433), .A4(n3499), 
        .ZN(n3317) );
  nr02d1 U4946 ( .A1(n3434), .A2(n3317), .ZN(n3255) );
  buffd1 U4947 ( .I(n3255), .Z(n3282) );
  nd02d1 U4948 ( .A1(n3499), .A2(n3251), .ZN(n3482) );
  buffd1 U4949 ( .I(n3482), .Z(n3500) );
  buffd1 U4950 ( .I(n3255), .Z(n3286) );
  aoim22d1 U4951 ( .A1(n3282), .A2(n3500), .B1(\RegFilePlugin_regFile[31][0] ), 
        .B2(n3286), .Z(n5228) );
  buffd1 U4952 ( .I(n3255), .Z(n3279) );
  nd02d1 U4953 ( .A1(n3499), .A2(n3252), .ZN(n3338) );
  aoim22d1 U4954 ( .A1(n3279), .A2(n3338), .B1(\RegFilePlugin_regFile[31][31] ), .B2(n3286), .Z(n5227) );
  nd02d1 U4955 ( .A1(n3499), .A2(n3253), .ZN(n3503) );
  aoim22d1 U4956 ( .A1(n3282), .A2(n3503), .B1(\RegFilePlugin_regFile[31][30] ), .B2(n3279), .Z(n5226) );
  nd02d1 U4957 ( .A1(n3499), .A2(n3254), .ZN(n3339) );
  buffd1 U4958 ( .I(n3339), .Z(n3505) );
  aoim22d1 U4959 ( .A1(n3282), .A2(n3505), .B1(\RegFilePlugin_regFile[31][29] ), .B2(n3279), .Z(n5225) );
  nd02d1 U4960 ( .A1(n3499), .A2(n3256), .ZN(n3476) );
  buffd1 U4961 ( .I(n3476), .Z(n3484) );
  aoim22d1 U4962 ( .A1(n3279), .A2(n3484), .B1(\RegFilePlugin_regFile[31][28] ), .B2(n3279), .Z(n5224) );
  nd02d1 U4963 ( .A1(n3499), .A2(n3257), .ZN(n3508) );
  aoim22d1 U4964 ( .A1(n3282), .A2(n3508), .B1(\RegFilePlugin_regFile[31][27] ), .B2(n3286), .Z(n5223) );
  nd02d1 U4965 ( .A1(n3499), .A2(n3258), .ZN(n3510) );
  aoim22d1 U4966 ( .A1(n3282), .A2(n3510), .B1(\RegFilePlugin_regFile[31][26] ), .B2(n3279), .Z(n5222) );
  nd02d1 U4967 ( .A1(n3499), .A2(n3259), .ZN(n3452) );
  buffd1 U4968 ( .I(n3452), .Z(n3512) );
  aoim22d1 U4969 ( .A1(n3279), .A2(n3512), .B1(\RegFilePlugin_regFile[31][25] ), .B2(n3255), .Z(n5221) );
  nd02d1 U4970 ( .A1(n3499), .A2(n3260), .ZN(n3341) );
  aoim22d1 U4971 ( .A1(n3279), .A2(n3341), .B1(\RegFilePlugin_regFile[31][24] ), .B2(n3282), .Z(n5220) );
  nd02d4 U4972 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3261), .ZN(n3454)
         );
  aoim22d1 U4973 ( .A1(n3282), .A2(n3454), .B1(\RegFilePlugin_regFile[31][23] ), .B2(n3255), .Z(n5219) );
  nd02d1 U4974 ( .A1(n3499), .A2(n3262), .ZN(n3455) );
  buffd1 U4975 ( .I(n3455), .Z(n3517) );
  aoim22d1 U4976 ( .A1(n3282), .A2(n3517), .B1(\RegFilePlugin_regFile[31][22] ), .B2(n3282), .Z(n5218) );
  buffd1 U4977 ( .I(n3342), .Z(n3519) );
  aoim22d1 U4978 ( .A1(n3282), .A2(n3519), .B1(\RegFilePlugin_regFile[31][21] ), .B2(n3282), .Z(n5217) );
  nd02d1 U4979 ( .A1(n3499), .A2(n3264), .ZN(n3343) );
  buffd1 U4980 ( .I(n3343), .Z(n3521) );
  aoim22d1 U4981 ( .A1(n3279), .A2(n3521), .B1(\RegFilePlugin_regFile[31][20] ), .B2(n3255), .Z(n5216) );
  buffd1 U4982 ( .I(n3344), .Z(n3523) );
  aoim22d1 U4983 ( .A1(n3255), .A2(n3523), .B1(\RegFilePlugin_regFile[31][19] ), .B2(n3282), .Z(n5215) );
  nd02d4 U4984 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3266), .ZN(n3456)
         );
  aoim22d1 U4985 ( .A1(n3286), .A2(n3456), .B1(\RegFilePlugin_regFile[31][18] ), .B2(n3282), .Z(n5214) );
  nd02d1 U4986 ( .A1(n3499), .A2(n3267), .ZN(n3457) );
  buffd1 U4987 ( .I(n3457), .Z(n3527) );
  aoim22d1 U4988 ( .A1(n3255), .A2(n3527), .B1(\RegFilePlugin_regFile[31][17] ), .B2(n3255), .Z(n5213) );
  buffd1 U4989 ( .I(n3458), .Z(n3529) );
  aoim22d1 U4990 ( .A1(n3282), .A2(n3529), .B1(\RegFilePlugin_regFile[31][16] ), .B2(n3255), .Z(n5212) );
  nd02d1 U4991 ( .A1(n3499), .A2(n3269), .ZN(n3366) );
  aoim22d1 U4992 ( .A1(n3279), .A2(n3366), .B1(\RegFilePlugin_regFile[31][15] ), .B2(n3255), .Z(n5211) );
  nd02d4 U4993 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3270), .ZN(n3459)
         );
  aoim22d1 U4994 ( .A1(n3255), .A2(n3459), .B1(\RegFilePlugin_regFile[31][14] ), .B2(n3255), .Z(n5210) );
  nd02d1 U4995 ( .A1(n3499), .A2(n3271), .ZN(n3485) );
  buffd1 U4996 ( .I(n3485), .Z(n3534) );
  aoim22d1 U4997 ( .A1(n3286), .A2(n3534), .B1(\RegFilePlugin_regFile[31][13] ), .B2(n3255), .Z(n5209) );
  nd02d4 U4998 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3272), .ZN(n3460)
         );
  aoim22d1 U4999 ( .A1(n3282), .A2(n3460), .B1(\RegFilePlugin_regFile[31][12] ), .B2(n3282), .Z(n5208) );
  nd02d4 U5000 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3273), .ZN(n3461)
         );
  aoim22d1 U5001 ( .A1(n3286), .A2(n3461), .B1(\RegFilePlugin_regFile[31][11] ), .B2(n3279), .Z(n5207) );
  nd02d4 U5002 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3274), .ZN(n3462)
         );
  aoim22d1 U5003 ( .A1(n3286), .A2(n3462), .B1(\RegFilePlugin_regFile[31][10] ), .B2(n3279), .Z(n5206) );
  nd02d4 U5004 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3275), .ZN(n3463)
         );
  aoim22d1 U5005 ( .A1(n3279), .A2(n3463), .B1(\RegFilePlugin_regFile[31][9] ), 
        .B2(n3279), .Z(n5205) );
  nd02d1 U5006 ( .A1(n3499), .A2(n3276), .ZN(n3464) );
  buffd1 U5007 ( .I(n3464), .Z(n3541) );
  aoim22d1 U5008 ( .A1(n3286), .A2(n3541), .B1(\RegFilePlugin_regFile[31][8] ), 
        .B2(n3279), .Z(n5204) );
  buffd1 U5009 ( .I(n3465), .Z(n3543) );
  aoim22d1 U5010 ( .A1(n3255), .A2(n3543), .B1(\RegFilePlugin_regFile[31][7] ), 
        .B2(n3279), .Z(n5203) );
  nd02d4 U5011 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3278), .ZN(n3467)
         );
  aoim22d1 U5012 ( .A1(n3286), .A2(n3467), .B1(\RegFilePlugin_regFile[31][6] ), 
        .B2(n3279), .Z(n5202) );
  nd02d4 U5013 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3280), .ZN(n3468)
         );
  aoim22d1 U5014 ( .A1(n3286), .A2(n3468), .B1(\RegFilePlugin_regFile[31][5] ), 
        .B2(n3286), .Z(n5201) );
  nd02d4 U5015 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3281), .ZN(n3469)
         );
  aoim22d1 U5016 ( .A1(n3282), .A2(n3469), .B1(\RegFilePlugin_regFile[31][4] ), 
        .B2(n3286), .Z(n5200) );
  nd02d1 U5017 ( .A1(n3499), .A2(n3283), .ZN(n3471) );
  buffd1 U5018 ( .I(n3471), .Z(n3551) );
  aoim22d1 U5019 ( .A1(n3255), .A2(n3551), .B1(\RegFilePlugin_regFile[31][3] ), 
        .B2(n3286), .Z(n5199) );
  nd02d4 U5020 ( .A1(IBusCachedPlugin_fetchPc_booted), .A2(n3284), .ZN(n3472)
         );
  aoim22d1 U5021 ( .A1(n3286), .A2(n3472), .B1(\RegFilePlugin_regFile[31][2] ), 
        .B2(n3286), .Z(n5198) );
  buffd1 U5022 ( .I(n3473), .Z(n3554) );
  aoim22d1 U5023 ( .A1(n3286), .A2(n3554), .B1(\RegFilePlugin_regFile[31][1] ), 
        .B2(n3286), .Z(n5197) );
  nr02d0 U5024 ( .A1(_zz_lastStageRegFileWrite_payload_address[7]), .A2(n3287), 
        .ZN(n3391) );
  nd03d0 U5025 ( .A1(_zz_lastStageRegFileWrite_payload_address[9]), .A2(
        _zz_lastStageRegFileWrite_payload_address[8]), .A3(n3391), .ZN(n3439)
         );
  nr02d1 U5026 ( .A1(n3317), .A2(n3439), .ZN(n3288) );
  buffd1 U5027 ( .I(n3288), .Z(n3289) );
  buffd1 U5028 ( .I(n3288), .Z(n3291) );
  aoim22d1 U5029 ( .A1(n3289), .A2(n3500), .B1(\RegFilePlugin_regFile[30][0] ), 
        .B2(n3291), .Z(n5196) );
  buffd1 U5030 ( .I(n3338), .Z(n3450) );
  aoim22d1 U5031 ( .A1(n3288), .A2(n3450), .B1(\RegFilePlugin_regFile[30][31] ), .B2(n3291), .Z(n5195) );
  buffd1 U5032 ( .I(n3503), .Z(n3490) );
  aoim22d1 U5033 ( .A1(n3289), .A2(n3490), .B1(\RegFilePlugin_regFile[30][30] ), .B2(n3288), .Z(n5194) );
  aoim22d1 U5034 ( .A1(n3289), .A2(n3505), .B1(\RegFilePlugin_regFile[30][29] ), .B2(n3288), .Z(n5193) );
  buffd1 U5035 ( .I(n3288), .Z(n3290) );
  aoim22d1 U5036 ( .A1(n3290), .A2(n3484), .B1(\RegFilePlugin_regFile[30][28] ), .B2(n3289), .Z(n5192) );
  buffd1 U5037 ( .I(n3508), .Z(n3492) );
  aoim22d1 U5038 ( .A1(n3289), .A2(n3492), .B1(\RegFilePlugin_regFile[30][27] ), .B2(n3290), .Z(n5191) );
  buffd1 U5039 ( .I(n3510), .Z(n3493) );
  aoim22d1 U5040 ( .A1(n3289), .A2(n3493), .B1(\RegFilePlugin_regFile[30][26] ), .B2(n3288), .Z(n5190) );
  aoim22d1 U5041 ( .A1(n3291), .A2(n3512), .B1(\RegFilePlugin_regFile[30][25] ), .B2(n3290), .Z(n5189) );
  buffd1 U5042 ( .I(n3341), .Z(n3453) );
  aoim22d1 U5043 ( .A1(n3288), .A2(n3453), .B1(\RegFilePlugin_regFile[30][24] ), .B2(n3289), .Z(n5188) );
  aoim22d1 U5044 ( .A1(n3289), .A2(n3454), .B1(\RegFilePlugin_regFile[30][23] ), .B2(n3290), .Z(n5187) );
  aoim22d1 U5045 ( .A1(n3289), .A2(n3517), .B1(\RegFilePlugin_regFile[30][22] ), .B2(n3289), .Z(n5186) );
  aoim22d1 U5046 ( .A1(n3289), .A2(n3342), .B1(\RegFilePlugin_regFile[30][21] ), .B2(n3289), .Z(n5185) );
  aoim22d1 U5047 ( .A1(n3288), .A2(n3343), .B1(\RegFilePlugin_regFile[30][20] ), .B2(n3290), .Z(n5184) );
  aoim22d1 U5048 ( .A1(n3290), .A2(n3344), .B1(\RegFilePlugin_regFile[30][19] ), .B2(n3289), .Z(n5183) );
  aoim22d1 U5049 ( .A1(n3291), .A2(n3456), .B1(\RegFilePlugin_regFile[30][18] ), .B2(n3289), .Z(n5182) );
  aoim22d1 U5050 ( .A1(n3290), .A2(n3527), .B1(\RegFilePlugin_regFile[30][17] ), .B2(n3290), .Z(n5181) );
  aoim22d1 U5051 ( .A1(n3289), .A2(n3458), .B1(\RegFilePlugin_regFile[30][16] ), .B2(n3290), .Z(n5180) );
  aoim22d1 U5052 ( .A1(n3288), .A2(n3366), .B1(\RegFilePlugin_regFile[30][15] ), .B2(n3290), .Z(n5179) );
  aoim22d1 U5053 ( .A1(n3290), .A2(n3459), .B1(\RegFilePlugin_regFile[30][14] ), .B2(n3290), .Z(n5178) );
  aoim22d1 U5054 ( .A1(n3291), .A2(n3534), .B1(\RegFilePlugin_regFile[30][13] ), .B2(n3290), .Z(n5177) );
  aoim22d1 U5055 ( .A1(n3289), .A2(n3460), .B1(\RegFilePlugin_regFile[30][12] ), .B2(n3290), .Z(n5176) );
  aoim22d1 U5056 ( .A1(n3291), .A2(n3461), .B1(\RegFilePlugin_regFile[30][11] ), .B2(n3288), .Z(n5175) );
  aoim22d1 U5057 ( .A1(n3291), .A2(n3462), .B1(\RegFilePlugin_regFile[30][10] ), .B2(n3288), .Z(n5174) );
  aoim22d1 U5058 ( .A1(n3288), .A2(n3463), .B1(\RegFilePlugin_regFile[30][9] ), 
        .B2(n3288), .Z(n5173) );
  aoim22d1 U5059 ( .A1(n3291), .A2(n3464), .B1(\RegFilePlugin_regFile[30][8] ), 
        .B2(n3290), .Z(n5172) );
  aoim22d1 U5060 ( .A1(n3290), .A2(n3465), .B1(\RegFilePlugin_regFile[30][7] ), 
        .B2(n3288), .Z(n5171) );
  aoim22d1 U5061 ( .A1(n3291), .A2(n3467), .B1(\RegFilePlugin_regFile[30][6] ), 
        .B2(n3288), .Z(n5170) );
  aoim22d1 U5062 ( .A1(n3291), .A2(n3468), .B1(\RegFilePlugin_regFile[30][5] ), 
        .B2(n3291), .Z(n5169) );
  aoim22d1 U5063 ( .A1(n3289), .A2(n3469), .B1(\RegFilePlugin_regFile[30][4] ), 
        .B2(n3291), .Z(n5168) );
  aoim22d1 U5064 ( .A1(n3290), .A2(n3471), .B1(\RegFilePlugin_regFile[30][3] ), 
        .B2(n3291), .Z(n5167) );
  aoim22d1 U5065 ( .A1(n3291), .A2(n3472), .B1(\RegFilePlugin_regFile[30][2] ), 
        .B2(n3291), .Z(n5166) );
  aoim22d1 U5066 ( .A1(n3291), .A2(n3473), .B1(\RegFilePlugin_regFile[30][1] ), 
        .B2(n3291), .Z(n5165) );
  inv0d0 U5067 ( .I(_zz_lastStageRegFileWrite_payload_address[8]), .ZN(n3314)
         );
  nd03d0 U5068 ( .A1(_zz_lastStageRegFileWrite_payload_address[9]), .A2(n3309), 
        .A3(n3314), .ZN(n3444) );
  nr02d1 U5069 ( .A1(n3317), .A2(n3444), .ZN(n3292) );
  buffd1 U5070 ( .I(n3292), .Z(n3293) );
  buffd1 U5071 ( .I(n3292), .Z(n3295) );
  aoim22d1 U5072 ( .A1(n3293), .A2(n3482), .B1(\RegFilePlugin_regFile[29][0] ), 
        .B2(n3295), .Z(n5164) );
  aoim22d1 U5073 ( .A1(n3292), .A2(n3338), .B1(\RegFilePlugin_regFile[29][31] ), .B2(n3295), .Z(n5163) );
  aoim22d1 U5074 ( .A1(n3293), .A2(n3503), .B1(\RegFilePlugin_regFile[29][30] ), .B2(n3293), .Z(n5162) );
  aoim22d1 U5075 ( .A1(n3293), .A2(n3505), .B1(\RegFilePlugin_regFile[29][29] ), .B2(n3292), .Z(n5161) );
  buffd1 U5076 ( .I(n3292), .Z(n3294) );
  aoim22d1 U5077 ( .A1(n3294), .A2(n3476), .B1(\RegFilePlugin_regFile[29][28] ), .B2(n3292), .Z(n5160) );
  aoim22d1 U5078 ( .A1(n3293), .A2(n3508), .B1(\RegFilePlugin_regFile[29][27] ), .B2(n3294), .Z(n5159) );
  aoim22d1 U5079 ( .A1(n3293), .A2(n3510), .B1(\RegFilePlugin_regFile[29][26] ), .B2(n3292), .Z(n5158) );
  aoim22d1 U5080 ( .A1(n3295), .A2(n3452), .B1(\RegFilePlugin_regFile[29][25] ), .B2(n3294), .Z(n5157) );
  aoim22d1 U5081 ( .A1(n3292), .A2(n3341), .B1(\RegFilePlugin_regFile[29][24] ), .B2(n3293), .Z(n5156) );
  aoim22d1 U5082 ( .A1(n3293), .A2(n3454), .B1(\RegFilePlugin_regFile[29][23] ), .B2(n3294), .Z(n5155) );
  aoim22d1 U5083 ( .A1(n3293), .A2(n3455), .B1(\RegFilePlugin_regFile[29][22] ), .B2(n3293), .Z(n5154) );
  aoim22d1 U5084 ( .A1(n3293), .A2(n3519), .B1(\RegFilePlugin_regFile[29][21] ), .B2(n3293), .Z(n5153) );
  aoim22d1 U5085 ( .A1(n3292), .A2(n3521), .B1(\RegFilePlugin_regFile[29][20] ), .B2(n3294), .Z(n5152) );
  aoim22d1 U5086 ( .A1(n3294), .A2(n3523), .B1(\RegFilePlugin_regFile[29][19] ), .B2(n3293), .Z(n5151) );
  aoim22d1 U5087 ( .A1(n3295), .A2(n3456), .B1(\RegFilePlugin_regFile[29][18] ), .B2(n3293), .Z(n5150) );
  aoim22d1 U5088 ( .A1(n3294), .A2(n3457), .B1(\RegFilePlugin_regFile[29][17] ), .B2(n3294), .Z(n5149) );
  aoim22d1 U5089 ( .A1(n3293), .A2(n3529), .B1(\RegFilePlugin_regFile[29][16] ), .B2(n3294), .Z(n5148) );
  aoim22d1 U5090 ( .A1(n3292), .A2(n3366), .B1(\RegFilePlugin_regFile[29][15] ), .B2(n3294), .Z(n5147) );
  aoim22d1 U5091 ( .A1(n3294), .A2(n3459), .B1(\RegFilePlugin_regFile[29][14] ), .B2(n3294), .Z(n5146) );
  aoim22d1 U5092 ( .A1(n3295), .A2(n3485), .B1(\RegFilePlugin_regFile[29][13] ), .B2(n3294), .Z(n5145) );
  aoim22d1 U5093 ( .A1(n3293), .A2(n3460), .B1(\RegFilePlugin_regFile[29][12] ), .B2(n3294), .Z(n5144) );
  aoim22d1 U5094 ( .A1(n3295), .A2(n3461), .B1(\RegFilePlugin_regFile[29][11] ), .B2(n3294), .Z(n5143) );
  aoim22d1 U5095 ( .A1(n3295), .A2(n3462), .B1(\RegFilePlugin_regFile[29][10] ), .B2(n3292), .Z(n5142) );
  aoim22d1 U5096 ( .A1(n3292), .A2(n3463), .B1(\RegFilePlugin_regFile[29][9] ), 
        .B2(n3292), .Z(n5141) );
  aoim22d1 U5097 ( .A1(n3295), .A2(n3541), .B1(\RegFilePlugin_regFile[29][8] ), 
        .B2(n3292), .Z(n5140) );
  aoim22d1 U5098 ( .A1(n3294), .A2(n3543), .B1(\RegFilePlugin_regFile[29][7] ), 
        .B2(n3292), .Z(n5139) );
  aoim22d1 U5099 ( .A1(n3295), .A2(n3467), .B1(\RegFilePlugin_regFile[29][6] ), 
        .B2(n3292), .Z(n5138) );
  aoim22d1 U5100 ( .A1(n3295), .A2(n3468), .B1(\RegFilePlugin_regFile[29][5] ), 
        .B2(n3295), .Z(n5137) );
  aoim22d1 U5101 ( .A1(n3293), .A2(n3469), .B1(\RegFilePlugin_regFile[29][4] ), 
        .B2(n3295), .Z(n5136) );
  aoim22d1 U5102 ( .A1(n3294), .A2(n3551), .B1(\RegFilePlugin_regFile[29][3] ), 
        .B2(n3295), .Z(n5135) );
  aoim22d1 U5103 ( .A1(n3295), .A2(n3472), .B1(\RegFilePlugin_regFile[29][2] ), 
        .B2(n3295), .Z(n5134) );
  aoim22d1 U5104 ( .A1(n3295), .A2(n3554), .B1(\RegFilePlugin_regFile[29][1] ), 
        .B2(n3295), .Z(n5133) );
  nd03d0 U5105 ( .A1(_zz_lastStageRegFileWrite_payload_address[9]), .A2(n3391), 
        .A3(n3314), .ZN(n3449) );
  buffd1 U5106 ( .I(n3296), .Z(n3298) );
  buffd1 U5107 ( .I(n3296), .Z(n3300) );
  aoim22d1 U5108 ( .A1(n3298), .A2(n3482), .B1(\RegFilePlugin_regFile[28][0] ), 
        .B2(n3300), .Z(n5132) );
  buffd1 U5109 ( .I(n3296), .Z(n3297) );
  aoim22d1 U5110 ( .A1(n3297), .A2(n3450), .B1(\RegFilePlugin_regFile[28][31] ), .B2(n3300), .Z(n5131) );
  aoim22d1 U5111 ( .A1(n3298), .A2(n3503), .B1(\RegFilePlugin_regFile[28][30] ), .B2(n3297), .Z(n5130) );
  aoim22d1 U5112 ( .A1(n3298), .A2(n3339), .B1(\RegFilePlugin_regFile[28][29] ), .B2(n3297), .Z(n5129) );
  buffd1 U5113 ( .I(n3296), .Z(n3299) );
  aoim22d1 U5114 ( .A1(n3299), .A2(n3476), .B1(\RegFilePlugin_regFile[28][28] ), .B2(n3297), .Z(n5128) );
  aoim22d1 U5115 ( .A1(n3298), .A2(n3508), .B1(\RegFilePlugin_regFile[28][27] ), .B2(n3299), .Z(n5127) );
  aoim22d1 U5116 ( .A1(n3298), .A2(n3510), .B1(\RegFilePlugin_regFile[28][26] ), .B2(n3297), .Z(n5126) );
  aoim22d1 U5117 ( .A1(n3297), .A2(n3512), .B1(\RegFilePlugin_regFile[28][25] ), .B2(n3299), .Z(n5125) );
  aoim22d1 U5118 ( .A1(n3297), .A2(n3453), .B1(\RegFilePlugin_regFile[28][24] ), .B2(n3298), .Z(n5124) );
  aoim22d1 U5119 ( .A1(n3298), .A2(n3454), .B1(\RegFilePlugin_regFile[28][23] ), .B2(n3299), .Z(n5123) );
  aoim22d1 U5120 ( .A1(n3298), .A2(n3517), .B1(\RegFilePlugin_regFile[28][22] ), .B2(n3298), .Z(n5122) );
  aoim22d1 U5121 ( .A1(n3298), .A2(n3342), .B1(\RegFilePlugin_regFile[28][21] ), .B2(n3298), .Z(n5121) );
  aoim22d1 U5122 ( .A1(n3297), .A2(n3521), .B1(\RegFilePlugin_regFile[28][20] ), .B2(n3299), .Z(n5120) );
  aoim22d1 U5123 ( .A1(n3299), .A2(n3344), .B1(\RegFilePlugin_regFile[28][19] ), .B2(n3298), .Z(n5119) );
  aoim22d1 U5124 ( .A1(n3300), .A2(n3456), .B1(\RegFilePlugin_regFile[28][18] ), .B2(n3298), .Z(n5118) );
  aoim22d1 U5125 ( .A1(n3299), .A2(n3527), .B1(\RegFilePlugin_regFile[28][17] ), .B2(n3299), .Z(n5117) );
  aoim22d1 U5126 ( .A1(n3298), .A2(n3458), .B1(\RegFilePlugin_regFile[28][16] ), .B2(n3299), .Z(n5116) );
  buffd1 U5127 ( .I(n3366), .Z(n3531) );
  aoim22d1 U5128 ( .A1(n3297), .A2(n3531), .B1(\RegFilePlugin_regFile[28][15] ), .B2(n3299), .Z(n5115) );
  aoim22d1 U5129 ( .A1(n3299), .A2(n3459), .B1(\RegFilePlugin_regFile[28][14] ), .B2(n3299), .Z(n5114) );
  aoim22d1 U5130 ( .A1(n3300), .A2(n3485), .B1(\RegFilePlugin_regFile[28][13] ), .B2(n3299), .Z(n5113) );
  aoim22d1 U5131 ( .A1(n3298), .A2(n3460), .B1(\RegFilePlugin_regFile[28][12] ), .B2(n3299), .Z(n5112) );
  aoim22d1 U5132 ( .A1(n3300), .A2(n3461), .B1(\RegFilePlugin_regFile[28][11] ), .B2(n3297), .Z(n5111) );
  aoim22d1 U5133 ( .A1(n3300), .A2(n3462), .B1(\RegFilePlugin_regFile[28][10] ), .B2(n3297), .Z(n5110) );
  aoim22d1 U5134 ( .A1(n3297), .A2(n3463), .B1(\RegFilePlugin_regFile[28][9] ), 
        .B2(n3297), .Z(n5109) );
  aoim22d1 U5135 ( .A1(n3300), .A2(n3464), .B1(\RegFilePlugin_regFile[28][8] ), 
        .B2(n3297), .Z(n5108) );
  aoim22d1 U5136 ( .A1(n3299), .A2(n3465), .B1(\RegFilePlugin_regFile[28][7] ), 
        .B2(n3297), .Z(n5107) );
  aoim22d1 U5137 ( .A1(n3300), .A2(n3467), .B1(\RegFilePlugin_regFile[28][6] ), 
        .B2(n3297), .Z(n5106) );
  aoim22d1 U5138 ( .A1(n3300), .A2(n3468), .B1(\RegFilePlugin_regFile[28][5] ), 
        .B2(n3300), .Z(n5105) );
  aoim22d1 U5139 ( .A1(n3298), .A2(n3469), .B1(\RegFilePlugin_regFile[28][4] ), 
        .B2(n3300), .Z(n5104) );
  aoim22d1 U5140 ( .A1(n3299), .A2(n3471), .B1(\RegFilePlugin_regFile[28][3] ), 
        .B2(n3300), .Z(n5103) );
  aoim22d1 U5141 ( .A1(n3300), .A2(n3472), .B1(\RegFilePlugin_regFile[28][2] ), 
        .B2(n3300), .Z(n5102) );
  aoim22d1 U5142 ( .A1(n3300), .A2(n3473), .B1(\RegFilePlugin_regFile[28][1] ), 
        .B2(n3300), .Z(n5101) );
  nd03d0 U5143 ( .A1(_zz_lastStageRegFileWrite_payload_address[8]), .A2(n3309), 
        .A3(n3315), .ZN(n3475) );
  nr02d1 U5144 ( .A1(n3317), .A2(n3475), .ZN(n3301) );
  buffd1 U5145 ( .I(n3301), .Z(n3303) );
  buffd1 U5146 ( .I(n3301), .Z(n3304) );
  aoim22d1 U5147 ( .A1(n3303), .A2(n3482), .B1(\RegFilePlugin_regFile[27][0] ), 
        .B2(n3304), .Z(n5100) );
  buffd1 U5148 ( .I(n3301), .Z(n3302) );
  aoim22d1 U5149 ( .A1(n3302), .A2(n3338), .B1(\RegFilePlugin_regFile[27][31] ), .B2(n3304), .Z(n5099) );
  aoim22d1 U5150 ( .A1(n3303), .A2(n3490), .B1(\RegFilePlugin_regFile[27][30] ), .B2(n3302), .Z(n5098) );
  aoim22d1 U5151 ( .A1(n3303), .A2(n3505), .B1(\RegFilePlugin_regFile[27][29] ), .B2(n3302), .Z(n5097) );
  aoim22d1 U5152 ( .A1(n3301), .A2(n3476), .B1(\RegFilePlugin_regFile[27][28] ), .B2(n3302), .Z(n5096) );
  aoim22d1 U5153 ( .A1(n3303), .A2(n3492), .B1(\RegFilePlugin_regFile[27][27] ), .B2(n3301), .Z(n5095) );
  aoim22d1 U5154 ( .A1(n3303), .A2(n3493), .B1(\RegFilePlugin_regFile[27][26] ), .B2(n3302), .Z(n5094) );
  aoim22d1 U5155 ( .A1(n3302), .A2(n3452), .B1(\RegFilePlugin_regFile[27][25] ), .B2(n3301), .Z(n5093) );
  aoim22d1 U5156 ( .A1(n3302), .A2(n3341), .B1(\RegFilePlugin_regFile[27][24] ), .B2(n3303), .Z(n5092) );
  aoim22d1 U5157 ( .A1(n3303), .A2(n3454), .B1(\RegFilePlugin_regFile[27][23] ), .B2(n3301), .Z(n5091) );
  aoim22d1 U5158 ( .A1(n3303), .A2(n3455), .B1(\RegFilePlugin_regFile[27][22] ), .B2(n3303), .Z(n5090) );
  aoim22d1 U5159 ( .A1(n3303), .A2(n3519), .B1(\RegFilePlugin_regFile[27][21] ), .B2(n3303), .Z(n5089) );
  aoim22d1 U5160 ( .A1(n3302), .A2(n3521), .B1(\RegFilePlugin_regFile[27][20] ), .B2(n3301), .Z(n5088) );
  aoim22d1 U5161 ( .A1(n3302), .A2(n3523), .B1(\RegFilePlugin_regFile[27][19] ), .B2(n3303), .Z(n5087) );
  aoim22d1 U5162 ( .A1(n3304), .A2(n3456), .B1(\RegFilePlugin_regFile[27][18] ), .B2(n3303), .Z(n5086) );
  aoim22d1 U5163 ( .A1(n3304), .A2(n3457), .B1(\RegFilePlugin_regFile[27][17] ), .B2(n3303), .Z(n5085) );
  aoim22d1 U5164 ( .A1(n3303), .A2(n3529), .B1(\RegFilePlugin_regFile[27][16] ), .B2(n3301), .Z(n5084) );
  aoim22d1 U5165 ( .A1(n3302), .A2(n3531), .B1(\RegFilePlugin_regFile[27][15] ), .B2(n3301), .Z(n5083) );
  aoim22d1 U5166 ( .A1(n3301), .A2(n3459), .B1(\RegFilePlugin_regFile[27][14] ), .B2(n3301), .Z(n5082) );
  aoim22d1 U5167 ( .A1(n3304), .A2(n3485), .B1(\RegFilePlugin_regFile[27][13] ), .B2(n3301), .Z(n5081) );
  aoim22d1 U5168 ( .A1(n3303), .A2(n3460), .B1(\RegFilePlugin_regFile[27][12] ), .B2(n3301), .Z(n5080) );
  aoim22d1 U5169 ( .A1(n3304), .A2(n3461), .B1(\RegFilePlugin_regFile[27][11] ), .B2(n3302), .Z(n5079) );
  aoim22d1 U5170 ( .A1(n3304), .A2(n3462), .B1(\RegFilePlugin_regFile[27][10] ), .B2(n3302), .Z(n5078) );
  aoim22d1 U5171 ( .A1(n3302), .A2(n3463), .B1(\RegFilePlugin_regFile[27][9] ), 
        .B2(n3302), .Z(n5077) );
  aoim22d1 U5172 ( .A1(n3304), .A2(n3541), .B1(\RegFilePlugin_regFile[27][8] ), 
        .B2(n3302), .Z(n5076) );
  aoim22d1 U5173 ( .A1(n3301), .A2(n3543), .B1(\RegFilePlugin_regFile[27][7] ), 
        .B2(n3302), .Z(n5075) );
  aoim22d1 U5174 ( .A1(n3304), .A2(n3467), .B1(\RegFilePlugin_regFile[27][6] ), 
        .B2(n3302), .Z(n5074) );
  aoim22d1 U5175 ( .A1(n3304), .A2(n3468), .B1(\RegFilePlugin_regFile[27][5] ), 
        .B2(n3304), .Z(n5073) );
  aoim22d1 U5176 ( .A1(n3303), .A2(n3469), .B1(\RegFilePlugin_regFile[27][4] ), 
        .B2(n3304), .Z(n5072) );
  aoim22d1 U5177 ( .A1(n3301), .A2(n3551), .B1(\RegFilePlugin_regFile[27][3] ), 
        .B2(n3304), .Z(n5071) );
  aoim22d1 U5178 ( .A1(n3304), .A2(n3472), .B1(\RegFilePlugin_regFile[27][2] ), 
        .B2(n3304), .Z(n5070) );
  aoim22d1 U5179 ( .A1(n3304), .A2(n3554), .B1(\RegFilePlugin_regFile[27][1] ), 
        .B2(n3304), .Z(n5069) );
  nd03d0 U5180 ( .A1(_zz_lastStageRegFileWrite_payload_address[8]), .A2(n3391), 
        .A3(n3315), .ZN(n3481) );
  nr02d1 U5181 ( .A1(n3317), .A2(n3481), .ZN(n3305) );
  buffd1 U5182 ( .I(n3305), .Z(n3307) );
  buffd1 U5183 ( .I(n3305), .Z(n3308) );
  aoim22d1 U5184 ( .A1(n3307), .A2(n3482), .B1(\RegFilePlugin_regFile[26][0] ), 
        .B2(n3308), .Z(n5068) );
  buffd1 U5185 ( .I(n3305), .Z(n3306) );
  aoim22d1 U5186 ( .A1(n3306), .A2(n3338), .B1(\RegFilePlugin_regFile[26][31] ), .B2(n3308), .Z(n5067) );
  aoim22d1 U5187 ( .A1(n3307), .A2(n3503), .B1(\RegFilePlugin_regFile[26][30] ), .B2(n3306), .Z(n5066) );
  aoim22d1 U5188 ( .A1(n3307), .A2(n3505), .B1(\RegFilePlugin_regFile[26][29] ), .B2(n3306), .Z(n5065) );
  aoim22d1 U5189 ( .A1(n3305), .A2(n3476), .B1(\RegFilePlugin_regFile[26][28] ), .B2(n3306), .Z(n5064) );
  aoim22d1 U5190 ( .A1(n3307), .A2(n3508), .B1(\RegFilePlugin_regFile[26][27] ), .B2(n3305), .Z(n5063) );
  aoim22d1 U5191 ( .A1(n3307), .A2(n3510), .B1(\RegFilePlugin_regFile[26][26] ), .B2(n3306), .Z(n5062) );
  aoim22d1 U5192 ( .A1(n3306), .A2(n3512), .B1(\RegFilePlugin_regFile[26][25] ), .B2(n3306), .Z(n5061) );
  aoim22d1 U5193 ( .A1(n3306), .A2(n3341), .B1(\RegFilePlugin_regFile[26][24] ), .B2(n3307), .Z(n5060) );
  aoim22d1 U5194 ( .A1(n3307), .A2(n3454), .B1(\RegFilePlugin_regFile[26][23] ), .B2(n3305), .Z(n5059) );
  aoim22d1 U5195 ( .A1(n3307), .A2(n3517), .B1(\RegFilePlugin_regFile[26][22] ), .B2(n3307), .Z(n5058) );
  aoim22d1 U5196 ( .A1(n3307), .A2(n3519), .B1(\RegFilePlugin_regFile[26][21] ), .B2(n3307), .Z(n5057) );
  aoim22d1 U5197 ( .A1(n3306), .A2(n3521), .B1(\RegFilePlugin_regFile[26][20] ), .B2(n3305), .Z(n5056) );
  aoim22d1 U5198 ( .A1(n3305), .A2(n3523), .B1(\RegFilePlugin_regFile[26][19] ), .B2(n3307), .Z(n5055) );
  aoim22d1 U5199 ( .A1(n3308), .A2(n3456), .B1(\RegFilePlugin_regFile[26][18] ), .B2(n3307), .Z(n5054) );
  aoim22d1 U5200 ( .A1(n3305), .A2(n3527), .B1(\RegFilePlugin_regFile[26][17] ), .B2(n3307), .Z(n5053) );
  aoim22d1 U5201 ( .A1(n3307), .A2(n3529), .B1(\RegFilePlugin_regFile[26][16] ), .B2(n3305), .Z(n5052) );
  aoim22d1 U5202 ( .A1(n3306), .A2(n3366), .B1(\RegFilePlugin_regFile[26][15] ), .B2(n3305), .Z(n5051) );
  aoim22d1 U5203 ( .A1(n3305), .A2(n3459), .B1(\RegFilePlugin_regFile[26][14] ), .B2(n3305), .Z(n5050) );
  aoim22d1 U5204 ( .A1(n3308), .A2(n3485), .B1(\RegFilePlugin_regFile[26][13] ), .B2(n3305), .Z(n5049) );
  aoim22d1 U5205 ( .A1(n3307), .A2(n3460), .B1(\RegFilePlugin_regFile[26][12] ), .B2(n3305), .Z(n5048) );
  aoim22d1 U5206 ( .A1(n3308), .A2(n3461), .B1(\RegFilePlugin_regFile[26][11] ), .B2(n3306), .Z(n5047) );
  aoim22d1 U5207 ( .A1(n3308), .A2(n3462), .B1(\RegFilePlugin_regFile[26][10] ), .B2(n3306), .Z(n5046) );
  aoim22d1 U5208 ( .A1(n3306), .A2(n3463), .B1(\RegFilePlugin_regFile[26][9] ), 
        .B2(n3306), .Z(n5045) );
  aoim22d1 U5209 ( .A1(n3308), .A2(n3541), .B1(\RegFilePlugin_regFile[26][8] ), 
        .B2(n3306), .Z(n5044) );
  aoim22d1 U5210 ( .A1(n3305), .A2(n3543), .B1(\RegFilePlugin_regFile[26][7] ), 
        .B2(n3306), .Z(n5043) );
  aoim22d1 U5211 ( .A1(n3308), .A2(n3467), .B1(\RegFilePlugin_regFile[26][6] ), 
        .B2(n3306), .Z(n5042) );
  aoim22d1 U5212 ( .A1(n3308), .A2(n3468), .B1(\RegFilePlugin_regFile[26][5] ), 
        .B2(n3308), .Z(n5041) );
  aoim22d1 U5213 ( .A1(n3307), .A2(n3469), .B1(\RegFilePlugin_regFile[26][4] ), 
        .B2(n3308), .Z(n5040) );
  aoim22d1 U5214 ( .A1(n3308), .A2(n3551), .B1(\RegFilePlugin_regFile[26][3] ), 
        .B2(n3308), .Z(n5039) );
  aoim22d1 U5215 ( .A1(n3308), .A2(n3472), .B1(\RegFilePlugin_regFile[26][2] ), 
        .B2(n3308), .Z(n5038) );
  aoim22d1 U5216 ( .A1(n3308), .A2(n3554), .B1(\RegFilePlugin_regFile[26][1] ), 
        .B2(n3308), .Z(n5037) );
  nr02d1 U5217 ( .A1(n3317), .A2(n3489), .ZN(n3310) );
  buffd1 U5218 ( .I(n3310), .Z(n3312) );
  aoim22d1 U5219 ( .A1(n3312), .A2(n3482), .B1(\RegFilePlugin_regFile[25][0] ), 
        .B2(n3310), .Z(n5036) );
  buffd1 U5220 ( .I(n3310), .Z(n3311) );
  aoim22d1 U5221 ( .A1(n3311), .A2(n3450), .B1(\RegFilePlugin_regFile[25][31] ), .B2(n3310), .Z(n5035) );
  aoim22d1 U5222 ( .A1(n3312), .A2(n3490), .B1(\RegFilePlugin_regFile[25][30] ), .B2(n3311), .Z(n5034) );
  aoim22d1 U5223 ( .A1(n3312), .A2(n3505), .B1(\RegFilePlugin_regFile[25][29] ), .B2(n3311), .Z(n5033) );
  buffd1 U5224 ( .I(n3310), .Z(n3313) );
  aoim22d1 U5225 ( .A1(n3313), .A2(n3476), .B1(\RegFilePlugin_regFile[25][28] ), .B2(n3311), .Z(n5032) );
  aoim22d1 U5226 ( .A1(n3312), .A2(n3492), .B1(\RegFilePlugin_regFile[25][27] ), .B2(n3313), .Z(n5031) );
  aoim22d1 U5227 ( .A1(n3312), .A2(n3493), .B1(\RegFilePlugin_regFile[25][26] ), .B2(n3311), .Z(n5030) );
  aoim22d1 U5228 ( .A1(n3311), .A2(n3452), .B1(\RegFilePlugin_regFile[25][25] ), .B2(n3313), .Z(n5029) );
  aoim22d1 U5229 ( .A1(n3311), .A2(n3453), .B1(\RegFilePlugin_regFile[25][24] ), .B2(n3312), .Z(n5028) );
  aoim22d1 U5230 ( .A1(n3312), .A2(n3454), .B1(\RegFilePlugin_regFile[25][23] ), .B2(n3313), .Z(n5027) );
  aoim22d1 U5231 ( .A1(n3312), .A2(n3455), .B1(\RegFilePlugin_regFile[25][22] ), .B2(n3312), .Z(n5026) );
  aoim22d1 U5232 ( .A1(n3312), .A2(n3342), .B1(\RegFilePlugin_regFile[25][21] ), .B2(n3312), .Z(n5025) );
  aoim22d1 U5233 ( .A1(n3311), .A2(n3343), .B1(\RegFilePlugin_regFile[25][20] ), .B2(n3313), .Z(n5024) );
  aoim22d1 U5234 ( .A1(n3313), .A2(n3344), .B1(\RegFilePlugin_regFile[25][19] ), .B2(n3312), .Z(n5023) );
  aoim22d1 U5235 ( .A1(n3310), .A2(n3456), .B1(\RegFilePlugin_regFile[25][18] ), .B2(n3312), .Z(n5022) );
  aoim22d1 U5236 ( .A1(n3313), .A2(n3457), .B1(\RegFilePlugin_regFile[25][17] ), .B2(n3313), .Z(n5021) );
  aoim22d1 U5237 ( .A1(n3312), .A2(n3529), .B1(\RegFilePlugin_regFile[25][16] ), .B2(n3313), .Z(n5020) );
  aoim22d1 U5238 ( .A1(n3311), .A2(n3531), .B1(\RegFilePlugin_regFile[25][15] ), .B2(n3313), .Z(n5019) );
  aoim22d1 U5239 ( .A1(n3313), .A2(n3459), .B1(\RegFilePlugin_regFile[25][14] ), .B2(n3313), .Z(n5018) );
  aoim22d1 U5240 ( .A1(n3310), .A2(n3485), .B1(\RegFilePlugin_regFile[25][13] ), .B2(n3313), .Z(n5017) );
  aoim22d1 U5241 ( .A1(n3312), .A2(n3460), .B1(\RegFilePlugin_regFile[25][12] ), .B2(n3313), .Z(n5016) );
  aoim22d1 U5242 ( .A1(n3313), .A2(n3461), .B1(\RegFilePlugin_regFile[25][11] ), .B2(n3311), .Z(n5015) );
  aoim22d1 U5243 ( .A1(n3310), .A2(n3462), .B1(\RegFilePlugin_regFile[25][10] ), .B2(n3311), .Z(n5014) );
  aoim22d1 U5244 ( .A1(n3311), .A2(n3463), .B1(\RegFilePlugin_regFile[25][9] ), 
        .B2(n3311), .Z(n5013) );
  aoim22d1 U5245 ( .A1(n3310), .A2(n3541), .B1(\RegFilePlugin_regFile[25][8] ), 
        .B2(n3311), .Z(n5012) );
  aoim22d1 U5246 ( .A1(n3313), .A2(n3543), .B1(\RegFilePlugin_regFile[25][7] ), 
        .B2(n3311), .Z(n5011) );
  aoim22d1 U5247 ( .A1(n3310), .A2(n3467), .B1(\RegFilePlugin_regFile[25][6] ), 
        .B2(n3311), .Z(n5010) );
  aoim22d1 U5248 ( .A1(n3310), .A2(n3468), .B1(\RegFilePlugin_regFile[25][5] ), 
        .B2(n3312), .Z(n5009) );
  aoim22d1 U5249 ( .A1(n3312), .A2(n3469), .B1(\RegFilePlugin_regFile[25][4] ), 
        .B2(n3311), .Z(n5008) );
  aoim22d1 U5250 ( .A1(n3313), .A2(n3551), .B1(\RegFilePlugin_regFile[25][3] ), 
        .B2(n3310), .Z(n5007) );
  aoim22d1 U5251 ( .A1(n3310), .A2(n3472), .B1(\RegFilePlugin_regFile[25][2] ), 
        .B2(n3310), .Z(n5006) );
  aoim22d1 U5252 ( .A1(n3310), .A2(n3554), .B1(\RegFilePlugin_regFile[25][1] ), 
        .B2(n3310), .Z(n5005) );
  nr02d1 U5253 ( .A1(n3317), .A2(n3498), .ZN(n3318) );
  buffd1 U5254 ( .I(n3318), .Z(n3320) );
  buffd1 U5255 ( .I(n3318), .Z(n3321) );
  aoim22d1 U5256 ( .A1(n3320), .A2(n3482), .B1(\RegFilePlugin_regFile[24][0] ), 
        .B2(n3321), .Z(n5004) );
  buffd1 U5257 ( .I(n3318), .Z(n3319) );
  aoim22d1 U5258 ( .A1(n3319), .A2(n3338), .B1(\RegFilePlugin_regFile[24][31] ), .B2(n3321), .Z(n5003) );
  aoim22d1 U5259 ( .A1(n3320), .A2(n3503), .B1(\RegFilePlugin_regFile[24][30] ), .B2(n3319), .Z(n5002) );
  aoim22d1 U5260 ( .A1(n3320), .A2(n3505), .B1(\RegFilePlugin_regFile[24][29] ), .B2(n3319), .Z(n5001) );
  aoim22d1 U5261 ( .A1(n3318), .A2(n3476), .B1(\RegFilePlugin_regFile[24][28] ), .B2(n3319), .Z(n5000) );
  aoim22d1 U5262 ( .A1(n3320), .A2(n3508), .B1(\RegFilePlugin_regFile[24][27] ), .B2(n3318), .Z(n4999) );
  aoim22d1 U5263 ( .A1(n3320), .A2(n3510), .B1(\RegFilePlugin_regFile[24][26] ), .B2(n3319), .Z(n4998) );
  aoim22d1 U5264 ( .A1(n3319), .A2(n3512), .B1(\RegFilePlugin_regFile[24][25] ), .B2(n3319), .Z(n4997) );
  aoim22d1 U5265 ( .A1(n3319), .A2(n3341), .B1(\RegFilePlugin_regFile[24][24] ), .B2(n3320), .Z(n4996) );
  aoim22d1 U5266 ( .A1(n3320), .A2(n3454), .B1(\RegFilePlugin_regFile[24][23] ), .B2(n3318), .Z(n4995) );
  aoim22d1 U5267 ( .A1(n3320), .A2(n3517), .B1(\RegFilePlugin_regFile[24][22] ), .B2(n3320), .Z(n4994) );
  aoim22d1 U5268 ( .A1(n3320), .A2(n3519), .B1(\RegFilePlugin_regFile[24][21] ), .B2(n3320), .Z(n4993) );
  aoim22d1 U5269 ( .A1(n3319), .A2(n3521), .B1(\RegFilePlugin_regFile[24][20] ), .B2(n3318), .Z(n4992) );
  aoim22d1 U5270 ( .A1(n3321), .A2(n3523), .B1(\RegFilePlugin_regFile[24][19] ), .B2(n3320), .Z(n4991) );
  aoim22d1 U5271 ( .A1(n3321), .A2(n3456), .B1(\RegFilePlugin_regFile[24][18] ), .B2(n3320), .Z(n4990) );
  aoim22d1 U5272 ( .A1(n3318), .A2(n3527), .B1(\RegFilePlugin_regFile[24][17] ), .B2(n3320), .Z(n4989) );
  aoim22d1 U5273 ( .A1(n3320), .A2(n3529), .B1(\RegFilePlugin_regFile[24][16] ), .B2(n3318), .Z(n4988) );
  aoim22d1 U5274 ( .A1(n3319), .A2(n3366), .B1(\RegFilePlugin_regFile[24][15] ), .B2(n3318), .Z(n4987) );
  aoim22d1 U5275 ( .A1(n3318), .A2(n3459), .B1(\RegFilePlugin_regFile[24][14] ), .B2(n3318), .Z(n4986) );
  aoim22d1 U5276 ( .A1(n3321), .A2(n3485), .B1(\RegFilePlugin_regFile[24][13] ), .B2(n3318), .Z(n4985) );
  aoim22d1 U5277 ( .A1(n3320), .A2(n3460), .B1(\RegFilePlugin_regFile[24][12] ), .B2(n3318), .Z(n4984) );
  aoim22d1 U5278 ( .A1(n3321), .A2(n3461), .B1(\RegFilePlugin_regFile[24][11] ), .B2(n3319), .Z(n4983) );
  aoim22d1 U5279 ( .A1(n3321), .A2(n3462), .B1(\RegFilePlugin_regFile[24][10] ), .B2(n3319), .Z(n4982) );
  aoim22d1 U5280 ( .A1(n3319), .A2(n3463), .B1(\RegFilePlugin_regFile[24][9] ), 
        .B2(n3319), .Z(n4981) );
  aoim22d1 U5281 ( .A1(n3321), .A2(n3541), .B1(\RegFilePlugin_regFile[24][8] ), 
        .B2(n3319), .Z(n4980) );
  aoim22d1 U5282 ( .A1(n3318), .A2(n3543), .B1(\RegFilePlugin_regFile[24][7] ), 
        .B2(n3319), .Z(n4979) );
  aoim22d1 U5283 ( .A1(n3321), .A2(n3467), .B1(\RegFilePlugin_regFile[24][6] ), 
        .B2(n3319), .Z(n4978) );
  aoim22d1 U5284 ( .A1(n3321), .A2(n3468), .B1(\RegFilePlugin_regFile[24][5] ), 
        .B2(n3321), .Z(n4977) );
  aoim22d1 U5285 ( .A1(n3320), .A2(n3469), .B1(\RegFilePlugin_regFile[24][4] ), 
        .B2(n3321), .Z(n4976) );
  aoim22d1 U5286 ( .A1(n3318), .A2(n3551), .B1(\RegFilePlugin_regFile[24][3] ), 
        .B2(n3321), .Z(n4975) );
  aoim22d1 U5287 ( .A1(n3321), .A2(n3472), .B1(\RegFilePlugin_regFile[24][2] ), 
        .B2(n3321), .Z(n4974) );
  aoim22d1 U5288 ( .A1(n3321), .A2(n3554), .B1(\RegFilePlugin_regFile[24][1] ), 
        .B2(n3321), .Z(n4973) );
  inv0d0 U5289 ( .I(_zz_lastStageRegFileWrite_payload_address[10]), .ZN(n3432)
         );
  nd04d0 U5290 ( .A1(_zz_lastStageRegFileWrite_payload_address[11]), .A2(n3433), .A3(n3499), .A4(n3432), .ZN(n3356) );
  nr02d1 U5291 ( .A1(n3434), .A2(n3356), .ZN(n3322) );
  buffd1 U5292 ( .I(n3322), .Z(n3324) );
  buffd1 U5293 ( .I(n3322), .Z(n3325) );
  aoim22d1 U5294 ( .A1(n3324), .A2(n3500), .B1(\RegFilePlugin_regFile[23][0] ), 
        .B2(n3325), .Z(n4972) );
  buffd1 U5295 ( .I(n3322), .Z(n3323) );
  aoim22d1 U5296 ( .A1(n3323), .A2(n3450), .B1(\RegFilePlugin_regFile[23][31] ), .B2(n3325), .Z(n4971) );
  aoim22d1 U5297 ( .A1(n3324), .A2(n3490), .B1(\RegFilePlugin_regFile[23][30] ), .B2(n3323), .Z(n4970) );
  aoim22d1 U5298 ( .A1(n3324), .A2(n3339), .B1(\RegFilePlugin_regFile[23][29] ), .B2(n3323), .Z(n4969) );
  aoim22d1 U5299 ( .A1(n3322), .A2(n3484), .B1(\RegFilePlugin_regFile[23][28] ), .B2(n3323), .Z(n4968) );
  aoim22d1 U5300 ( .A1(n3324), .A2(n3492), .B1(\RegFilePlugin_regFile[23][27] ), .B2(n3322), .Z(n4967) );
  aoim22d1 U5301 ( .A1(n3324), .A2(n3493), .B1(\RegFilePlugin_regFile[23][26] ), .B2(n3323), .Z(n4966) );
  aoim22d1 U5302 ( .A1(n3323), .A2(n3512), .B1(\RegFilePlugin_regFile[23][25] ), .B2(n3325), .Z(n4965) );
  aoim22d1 U5303 ( .A1(n3323), .A2(n3453), .B1(\RegFilePlugin_regFile[23][24] ), .B2(n3324), .Z(n4964) );
  aoim22d1 U5304 ( .A1(n3324), .A2(n3454), .B1(\RegFilePlugin_regFile[23][23] ), .B2(n3322), .Z(n4963) );
  aoim22d1 U5305 ( .A1(n3324), .A2(n3517), .B1(\RegFilePlugin_regFile[23][22] ), .B2(n3324), .Z(n4962) );
  aoim22d1 U5306 ( .A1(n3324), .A2(n3342), .B1(\RegFilePlugin_regFile[23][21] ), .B2(n3324), .Z(n4961) );
  aoim22d1 U5307 ( .A1(n3323), .A2(n3343), .B1(\RegFilePlugin_regFile[23][20] ), .B2(n3322), .Z(n4960) );
  aoim22d1 U5308 ( .A1(n3322), .A2(n3344), .B1(\RegFilePlugin_regFile[23][19] ), .B2(n3324), .Z(n4959) );
  aoim22d1 U5309 ( .A1(n3325), .A2(n3456), .B1(\RegFilePlugin_regFile[23][18] ), .B2(n3324), .Z(n4958) );
  aoim22d1 U5310 ( .A1(n3322), .A2(n3527), .B1(\RegFilePlugin_regFile[23][17] ), .B2(n3322), .Z(n4957) );
  aoim22d1 U5311 ( .A1(n3324), .A2(n3529), .B1(\RegFilePlugin_regFile[23][16] ), .B2(n3323), .Z(n4956) );
  aoim22d1 U5312 ( .A1(n3323), .A2(n3366), .B1(\RegFilePlugin_regFile[23][15] ), .B2(n3322), .Z(n4955) );
  aoim22d1 U5313 ( .A1(n3322), .A2(n3459), .B1(\RegFilePlugin_regFile[23][14] ), .B2(n3324), .Z(n4954) );
  aoim22d1 U5314 ( .A1(n3325), .A2(n3485), .B1(\RegFilePlugin_regFile[23][13] ), .B2(n3322), .Z(n4953) );
  aoim22d1 U5315 ( .A1(n3324), .A2(n3460), .B1(\RegFilePlugin_regFile[23][12] ), .B2(n3322), .Z(n4952) );
  aoim22d1 U5316 ( .A1(n3325), .A2(n3461), .B1(\RegFilePlugin_regFile[23][11] ), .B2(n3323), .Z(n4951) );
  aoim22d1 U5317 ( .A1(n3325), .A2(n3462), .B1(\RegFilePlugin_regFile[23][10] ), .B2(n3323), .Z(n4950) );
  aoim22d1 U5318 ( .A1(n3323), .A2(n3463), .B1(\RegFilePlugin_regFile[23][9] ), 
        .B2(n3323), .Z(n4949) );
  aoim22d1 U5319 ( .A1(n3325), .A2(n3541), .B1(\RegFilePlugin_regFile[23][8] ), 
        .B2(n3323), .Z(n4948) );
  aoim22d1 U5320 ( .A1(n3322), .A2(n3543), .B1(\RegFilePlugin_regFile[23][7] ), 
        .B2(n3323), .Z(n4947) );
  aoim22d1 U5321 ( .A1(n3325), .A2(n3467), .B1(\RegFilePlugin_regFile[23][6] ), 
        .B2(n3323), .Z(n4946) );
  aoim22d1 U5322 ( .A1(n3325), .A2(n3468), .B1(\RegFilePlugin_regFile[23][5] ), 
        .B2(n3325), .Z(n4945) );
  aoim22d1 U5323 ( .A1(n3324), .A2(n3469), .B1(\RegFilePlugin_regFile[23][4] ), 
        .B2(n3325), .Z(n4944) );
  aoim22d1 U5324 ( .A1(n3322), .A2(n3551), .B1(\RegFilePlugin_regFile[23][3] ), 
        .B2(n3325), .Z(n4943) );
  aoim22d1 U5325 ( .A1(n3325), .A2(n3472), .B1(\RegFilePlugin_regFile[23][2] ), 
        .B2(n3325), .Z(n4942) );
  aoim22d1 U5326 ( .A1(n3325), .A2(n3554), .B1(\RegFilePlugin_regFile[23][1] ), 
        .B2(n3325), .Z(n4941) );
  nr02d1 U5327 ( .A1(n3439), .A2(n3356), .ZN(n3326) );
  buffd1 U5328 ( .I(n3326), .Z(n3328) );
  buffd1 U5329 ( .I(n3326), .Z(n3329) );
  aoim22d1 U5330 ( .A1(n3328), .A2(n3500), .B1(\RegFilePlugin_regFile[22][0] ), 
        .B2(n3329), .Z(n4940) );
  buffd1 U5331 ( .I(n3326), .Z(n3327) );
  aoim22d1 U5332 ( .A1(n3327), .A2(n3338), .B1(\RegFilePlugin_regFile[22][31] ), .B2(n3329), .Z(n4939) );
  aoim22d1 U5333 ( .A1(n3328), .A2(n3503), .B1(\RegFilePlugin_regFile[22][30] ), .B2(n3327), .Z(n4938) );
  aoim22d1 U5334 ( .A1(n3328), .A2(n3339), .B1(\RegFilePlugin_regFile[22][29] ), .B2(n3327), .Z(n4937) );
  aoim22d1 U5335 ( .A1(n3326), .A2(n3484), .B1(\RegFilePlugin_regFile[22][28] ), .B2(n3327), .Z(n4936) );
  aoim22d1 U5336 ( .A1(n3328), .A2(n3508), .B1(\RegFilePlugin_regFile[22][27] ), .B2(n3326), .Z(n4935) );
  aoim22d1 U5337 ( .A1(n3328), .A2(n3510), .B1(\RegFilePlugin_regFile[22][26] ), .B2(n3327), .Z(n4934) );
  aoim22d1 U5338 ( .A1(n3327), .A2(n3452), .B1(\RegFilePlugin_regFile[22][25] ), .B2(n3326), .Z(n4933) );
  aoim22d1 U5339 ( .A1(n3327), .A2(n3341), .B1(\RegFilePlugin_regFile[22][24] ), .B2(n3328), .Z(n4932) );
  aoim22d1 U5340 ( .A1(n3328), .A2(n3454), .B1(\RegFilePlugin_regFile[22][23] ), .B2(n3326), .Z(n4931) );
  aoim22d1 U5341 ( .A1(n3328), .A2(n3455), .B1(\RegFilePlugin_regFile[22][22] ), .B2(n3328), .Z(n4930) );
  aoim22d1 U5342 ( .A1(n3328), .A2(n3342), .B1(\RegFilePlugin_regFile[22][21] ), .B2(n3328), .Z(n4929) );
  aoim22d1 U5343 ( .A1(n3327), .A2(n3343), .B1(\RegFilePlugin_regFile[22][20] ), .B2(n3326), .Z(n4928) );
  aoim22d1 U5344 ( .A1(n3327), .A2(n3344), .B1(\RegFilePlugin_regFile[22][19] ), .B2(n3328), .Z(n4927) );
  aoim22d1 U5345 ( .A1(n3329), .A2(n3456), .B1(\RegFilePlugin_regFile[22][18] ), .B2(n3328), .Z(n4926) );
  aoim22d1 U5346 ( .A1(n3329), .A2(n3457), .B1(\RegFilePlugin_regFile[22][17] ), .B2(n3328), .Z(n4925) );
  aoim22d1 U5347 ( .A1(n3328), .A2(n3529), .B1(\RegFilePlugin_regFile[22][16] ), .B2(n3326), .Z(n4924) );
  aoim22d1 U5348 ( .A1(n3327), .A2(n3366), .B1(\RegFilePlugin_regFile[22][15] ), .B2(n3326), .Z(n4923) );
  aoim22d1 U5349 ( .A1(n3326), .A2(n3459), .B1(\RegFilePlugin_regFile[22][14] ), .B2(n3326), .Z(n4922) );
  aoim22d1 U5350 ( .A1(n3329), .A2(n3485), .B1(\RegFilePlugin_regFile[22][13] ), .B2(n3326), .Z(n4921) );
  aoim22d1 U5351 ( .A1(n3328), .A2(n3460), .B1(\RegFilePlugin_regFile[22][12] ), .B2(n3326), .Z(n4920) );
  aoim22d1 U5352 ( .A1(n3329), .A2(n3461), .B1(\RegFilePlugin_regFile[22][11] ), .B2(n3327), .Z(n4919) );
  aoim22d1 U5353 ( .A1(n3329), .A2(n3462), .B1(\RegFilePlugin_regFile[22][10] ), .B2(n3327), .Z(n4918) );
  aoim22d1 U5354 ( .A1(n3327), .A2(n3463), .B1(\RegFilePlugin_regFile[22][9] ), 
        .B2(n3327), .Z(n4917) );
  aoim22d1 U5355 ( .A1(n3329), .A2(n3541), .B1(\RegFilePlugin_regFile[22][8] ), 
        .B2(n3327), .Z(n4916) );
  aoim22d1 U5356 ( .A1(n3326), .A2(n3543), .B1(\RegFilePlugin_regFile[22][7] ), 
        .B2(n3327), .Z(n4915) );
  aoim22d1 U5357 ( .A1(n3329), .A2(n3467), .B1(\RegFilePlugin_regFile[22][6] ), 
        .B2(n3327), .Z(n4914) );
  aoim22d1 U5358 ( .A1(n3329), .A2(n3468), .B1(\RegFilePlugin_regFile[22][5] ), 
        .B2(n3329), .Z(n4913) );
  aoim22d1 U5359 ( .A1(n3328), .A2(n3469), .B1(\RegFilePlugin_regFile[22][4] ), 
        .B2(n3329), .Z(n4912) );
  aoim22d1 U5360 ( .A1(n3326), .A2(n3551), .B1(\RegFilePlugin_regFile[22][3] ), 
        .B2(n3329), .Z(n4911) );
  aoim22d1 U5361 ( .A1(n3329), .A2(n3472), .B1(\RegFilePlugin_regFile[22][2] ), 
        .B2(n3329), .Z(n4910) );
  aoim22d1 U5362 ( .A1(n3329), .A2(n3554), .B1(\RegFilePlugin_regFile[22][1] ), 
        .B2(n3329), .Z(n4909) );
  nr02d1 U5363 ( .A1(n3444), .A2(n3356), .ZN(n3330) );
  buffd1 U5364 ( .I(n3330), .Z(n3332) );
  buffd1 U5365 ( .I(n3330), .Z(n3333) );
  aoim22d1 U5366 ( .A1(n3332), .A2(n3500), .B1(\RegFilePlugin_regFile[21][0] ), 
        .B2(n3333), .Z(n4908) );
  buffd1 U5367 ( .I(n3330), .Z(n3331) );
  aoim22d1 U5368 ( .A1(n3331), .A2(n3450), .B1(\RegFilePlugin_regFile[21][31] ), .B2(n3333), .Z(n4907) );
  aoim22d1 U5369 ( .A1(n3332), .A2(n3503), .B1(\RegFilePlugin_regFile[21][30] ), .B2(n3331), .Z(n4906) );
  aoim22d1 U5370 ( .A1(n3332), .A2(n3339), .B1(\RegFilePlugin_regFile[21][29] ), .B2(n3331), .Z(n4905) );
  aoim22d1 U5371 ( .A1(n3330), .A2(n3484), .B1(\RegFilePlugin_regFile[21][28] ), .B2(n3331), .Z(n4904) );
  aoim22d1 U5372 ( .A1(n3332), .A2(n3508), .B1(\RegFilePlugin_regFile[21][27] ), .B2(n3330), .Z(n4903) );
  aoim22d1 U5373 ( .A1(n3332), .A2(n3510), .B1(\RegFilePlugin_regFile[21][26] ), .B2(n3331), .Z(n4902) );
  aoim22d1 U5374 ( .A1(n3331), .A2(n3452), .B1(\RegFilePlugin_regFile[21][25] ), .B2(n3332), .Z(n4901) );
  aoim22d1 U5375 ( .A1(n3331), .A2(n3453), .B1(\RegFilePlugin_regFile[21][24] ), .B2(n3332), .Z(n4900) );
  aoim22d1 U5376 ( .A1(n3332), .A2(n3454), .B1(\RegFilePlugin_regFile[21][23] ), .B2(n3330), .Z(n4899) );
  aoim22d1 U5377 ( .A1(n3332), .A2(n3455), .B1(\RegFilePlugin_regFile[21][22] ), .B2(n3332), .Z(n4898) );
  aoim22d1 U5378 ( .A1(n3332), .A2(n3342), .B1(\RegFilePlugin_regFile[21][21] ), .B2(n3332), .Z(n4897) );
  aoim22d1 U5379 ( .A1(n3331), .A2(n3343), .B1(\RegFilePlugin_regFile[21][20] ), .B2(n3330), .Z(n4896) );
  aoim22d1 U5380 ( .A1(n3330), .A2(n3344), .B1(\RegFilePlugin_regFile[21][19] ), .B2(n3332), .Z(n4895) );
  aoim22d1 U5381 ( .A1(n3333), .A2(n3456), .B1(\RegFilePlugin_regFile[21][18] ), .B2(n3332), .Z(n4894) );
  aoim22d1 U5382 ( .A1(n3330), .A2(n3457), .B1(\RegFilePlugin_regFile[21][17] ), .B2(n3330), .Z(n4893) );
  aoim22d1 U5383 ( .A1(n3332), .A2(n3458), .B1(\RegFilePlugin_regFile[21][16] ), .B2(n3331), .Z(n4892) );
  aoim22d1 U5384 ( .A1(n3331), .A2(n3366), .B1(\RegFilePlugin_regFile[21][15] ), .B2(n3330), .Z(n4891) );
  aoim22d1 U5385 ( .A1(n3330), .A2(n3459), .B1(\RegFilePlugin_regFile[21][14] ), .B2(n3330), .Z(n4890) );
  aoim22d1 U5386 ( .A1(n3333), .A2(n3485), .B1(\RegFilePlugin_regFile[21][13] ), .B2(n3330), .Z(n4889) );
  aoim22d1 U5387 ( .A1(n3332), .A2(n3460), .B1(\RegFilePlugin_regFile[21][12] ), .B2(n3330), .Z(n4888) );
  aoim22d1 U5388 ( .A1(n3333), .A2(n3461), .B1(\RegFilePlugin_regFile[21][11] ), .B2(n3331), .Z(n4887) );
  aoim22d1 U5389 ( .A1(n3333), .A2(n3462), .B1(\RegFilePlugin_regFile[21][10] ), .B2(n3331), .Z(n4886) );
  aoim22d1 U5390 ( .A1(n3331), .A2(n3463), .B1(\RegFilePlugin_regFile[21][9] ), 
        .B2(n3331), .Z(n4885) );
  aoim22d1 U5391 ( .A1(n3333), .A2(n3464), .B1(\RegFilePlugin_regFile[21][8] ), 
        .B2(n3331), .Z(n4884) );
  aoim22d1 U5392 ( .A1(n3330), .A2(n3465), .B1(\RegFilePlugin_regFile[21][7] ), 
        .B2(n3331), .Z(n4883) );
  aoim22d1 U5393 ( .A1(n3333), .A2(n3467), .B1(\RegFilePlugin_regFile[21][6] ), 
        .B2(n3331), .Z(n4882) );
  aoim22d1 U5394 ( .A1(n3333), .A2(n3468), .B1(\RegFilePlugin_regFile[21][5] ), 
        .B2(n3333), .Z(n4881) );
  aoim22d1 U5395 ( .A1(n3332), .A2(n3469), .B1(\RegFilePlugin_regFile[21][4] ), 
        .B2(n3333), .Z(n4880) );
  aoim22d1 U5396 ( .A1(n3333), .A2(n3471), .B1(\RegFilePlugin_regFile[21][3] ), 
        .B2(n3333), .Z(n4879) );
  aoim22d1 U5397 ( .A1(n3333), .A2(n3472), .B1(\RegFilePlugin_regFile[21][2] ), 
        .B2(n3333), .Z(n4878) );
  aoim22d1 U5398 ( .A1(n3333), .A2(n3473), .B1(\RegFilePlugin_regFile[21][1] ), 
        .B2(n3333), .Z(n4877) );
  nr02d1 U5399 ( .A1(n3449), .A2(n3356), .ZN(n3334) );
  buffd1 U5400 ( .I(n3334), .Z(n3336) );
  buffd1 U5401 ( .I(n3334), .Z(n3337) );
  aoim22d1 U5402 ( .A1(n3336), .A2(n3500), .B1(\RegFilePlugin_regFile[20][0] ), 
        .B2(n3337), .Z(n4876) );
  buffd1 U5403 ( .I(n3334), .Z(n3335) );
  aoim22d1 U5404 ( .A1(n3335), .A2(n3450), .B1(\RegFilePlugin_regFile[20][31] ), .B2(n3337), .Z(n4875) );
  aoim22d1 U5405 ( .A1(n3336), .A2(n3503), .B1(\RegFilePlugin_regFile[20][30] ), .B2(n3335), .Z(n4874) );
  aoim22d1 U5406 ( .A1(n3336), .A2(n3505), .B1(\RegFilePlugin_regFile[20][29] ), .B2(n3335), .Z(n4873) );
  aoim22d1 U5407 ( .A1(n3334), .A2(n3484), .B1(\RegFilePlugin_regFile[20][28] ), .B2(n3335), .Z(n4872) );
  aoim22d1 U5408 ( .A1(n3336), .A2(n3508), .B1(\RegFilePlugin_regFile[20][27] ), .B2(n3334), .Z(n4871) );
  aoim22d1 U5409 ( .A1(n3336), .A2(n3510), .B1(\RegFilePlugin_regFile[20][26] ), .B2(n3335), .Z(n4870) );
  aoim22d1 U5410 ( .A1(n3335), .A2(n3512), .B1(\RegFilePlugin_regFile[20][25] ), .B2(n3336), .Z(n4869) );
  aoim22d1 U5411 ( .A1(n3335), .A2(n3341), .B1(\RegFilePlugin_regFile[20][24] ), .B2(n3336), .Z(n4868) );
  aoim22d1 U5412 ( .A1(n3336), .A2(n3454), .B1(\RegFilePlugin_regFile[20][23] ), .B2(n3334), .Z(n4867) );
  aoim22d1 U5413 ( .A1(n3336), .A2(n3517), .B1(\RegFilePlugin_regFile[20][22] ), .B2(n3336), .Z(n4866) );
  aoim22d1 U5414 ( .A1(n3336), .A2(n3519), .B1(\RegFilePlugin_regFile[20][21] ), .B2(n3336), .Z(n4865) );
  aoim22d1 U5415 ( .A1(n3335), .A2(n3521), .B1(\RegFilePlugin_regFile[20][20] ), .B2(n3334), .Z(n4864) );
  aoim22d1 U5416 ( .A1(n3334), .A2(n3523), .B1(\RegFilePlugin_regFile[20][19] ), .B2(n3336), .Z(n4863) );
  aoim22d1 U5417 ( .A1(n3337), .A2(n3456), .B1(\RegFilePlugin_regFile[20][18] ), .B2(n3336), .Z(n4862) );
  aoim22d1 U5418 ( .A1(n3334), .A2(n3527), .B1(\RegFilePlugin_regFile[20][17] ), .B2(n3334), .Z(n4861) );
  aoim22d1 U5419 ( .A1(n3336), .A2(n3458), .B1(\RegFilePlugin_regFile[20][16] ), .B2(n3337), .Z(n4860) );
  aoim22d1 U5420 ( .A1(n3335), .A2(n3366), .B1(\RegFilePlugin_regFile[20][15] ), .B2(n3334), .Z(n4859) );
  aoim22d1 U5421 ( .A1(n3334), .A2(n3459), .B1(\RegFilePlugin_regFile[20][14] ), .B2(n3334), .Z(n4858) );
  aoim22d1 U5422 ( .A1(n3337), .A2(n3485), .B1(\RegFilePlugin_regFile[20][13] ), .B2(n3335), .Z(n4857) );
  aoim22d1 U5423 ( .A1(n3336), .A2(n3460), .B1(\RegFilePlugin_regFile[20][12] ), .B2(n3334), .Z(n4856) );
  aoim22d1 U5424 ( .A1(n3337), .A2(n3461), .B1(\RegFilePlugin_regFile[20][11] ), .B2(n3335), .Z(n4855) );
  aoim22d1 U5425 ( .A1(n3337), .A2(n3462), .B1(\RegFilePlugin_regFile[20][10] ), .B2(n3335), .Z(n4854) );
  aoim22d1 U5426 ( .A1(n3335), .A2(n3463), .B1(\RegFilePlugin_regFile[20][9] ), 
        .B2(n3335), .Z(n4853) );
  aoim22d1 U5427 ( .A1(n3337), .A2(n3464), .B1(\RegFilePlugin_regFile[20][8] ), 
        .B2(n3335), .Z(n4852) );
  aoim22d1 U5428 ( .A1(n3334), .A2(n3465), .B1(\RegFilePlugin_regFile[20][7] ), 
        .B2(n3335), .Z(n4851) );
  aoim22d1 U5429 ( .A1(n3337), .A2(n3467), .B1(\RegFilePlugin_regFile[20][6] ), 
        .B2(n3335), .Z(n4850) );
  aoim22d1 U5430 ( .A1(n3337), .A2(n3468), .B1(\RegFilePlugin_regFile[20][5] ), 
        .B2(n3337), .Z(n4849) );
  aoim22d1 U5431 ( .A1(n3336), .A2(n3469), .B1(\RegFilePlugin_regFile[20][4] ), 
        .B2(n3337), .Z(n4848) );
  aoim22d1 U5432 ( .A1(n3334), .A2(n3471), .B1(\RegFilePlugin_regFile[20][3] ), 
        .B2(n3337), .Z(n4847) );
  aoim22d1 U5433 ( .A1(n3337), .A2(n3472), .B1(\RegFilePlugin_regFile[20][2] ), 
        .B2(n3337), .Z(n4846) );
  aoim22d1 U5434 ( .A1(n3337), .A2(n3473), .B1(\RegFilePlugin_regFile[20][1] ), 
        .B2(n3337), .Z(n4845) );
  nr02d1 U5435 ( .A1(n3475), .A2(n3356), .ZN(n3340) );
  buffd1 U5436 ( .I(n3340), .Z(n3346) );
  buffd1 U5437 ( .I(n3340), .Z(n3347) );
  aoim22d1 U5438 ( .A1(n3346), .A2(n3500), .B1(\RegFilePlugin_regFile[19][0] ), 
        .B2(n3347), .Z(n4844) );
  buffd1 U5439 ( .I(n3340), .Z(n3345) );
  aoim22d1 U5440 ( .A1(n3345), .A2(n3338), .B1(\RegFilePlugin_regFile[19][31] ), .B2(n3347), .Z(n4843) );
  aoim22d1 U5441 ( .A1(n3346), .A2(n3503), .B1(\RegFilePlugin_regFile[19][30] ), .B2(n3345), .Z(n4842) );
  aoim22d1 U5442 ( .A1(n3346), .A2(n3339), .B1(\RegFilePlugin_regFile[19][29] ), .B2(n3345), .Z(n4841) );
  aoim22d1 U5443 ( .A1(n3340), .A2(n3484), .B1(\RegFilePlugin_regFile[19][28] ), .B2(n3345), .Z(n4840) );
  aoim22d1 U5444 ( .A1(n3346), .A2(n3508), .B1(\RegFilePlugin_regFile[19][27] ), .B2(n3340), .Z(n4839) );
  aoim22d1 U5445 ( .A1(n3346), .A2(n3510), .B1(\RegFilePlugin_regFile[19][26] ), .B2(n3345), .Z(n4838) );
  aoim22d1 U5446 ( .A1(n3345), .A2(n3452), .B1(\RegFilePlugin_regFile[19][25] ), .B2(n3345), .Z(n4837) );
  aoim22d1 U5447 ( .A1(n3345), .A2(n3341), .B1(\RegFilePlugin_regFile[19][24] ), .B2(n3346), .Z(n4836) );
  aoim22d1 U5448 ( .A1(n3346), .A2(n3454), .B1(\RegFilePlugin_regFile[19][23] ), .B2(n3340), .Z(n4835) );
  aoim22d1 U5449 ( .A1(n3346), .A2(n3455), .B1(\RegFilePlugin_regFile[19][22] ), .B2(n3346), .Z(n4834) );
  aoim22d1 U5450 ( .A1(n3346), .A2(n3342), .B1(\RegFilePlugin_regFile[19][21] ), .B2(n3346), .Z(n4833) );
  aoim22d1 U5451 ( .A1(n3345), .A2(n3343), .B1(\RegFilePlugin_regFile[19][20] ), .B2(n3340), .Z(n4832) );
  aoim22d1 U5452 ( .A1(n3340), .A2(n3344), .B1(\RegFilePlugin_regFile[19][19] ), .B2(n3346), .Z(n4831) );
  aoim22d1 U5453 ( .A1(n3347), .A2(n3456), .B1(\RegFilePlugin_regFile[19][18] ), .B2(n3346), .Z(n4830) );
  aoim22d1 U5454 ( .A1(n3340), .A2(n3457), .B1(\RegFilePlugin_regFile[19][17] ), .B2(n3340), .Z(n4829) );
  aoim22d1 U5455 ( .A1(n3346), .A2(n3529), .B1(\RegFilePlugin_regFile[19][16] ), .B2(n3347), .Z(n4828) );
  aoim22d1 U5456 ( .A1(n3345), .A2(n3366), .B1(\RegFilePlugin_regFile[19][15] ), .B2(n3340), .Z(n4827) );
  aoim22d1 U5457 ( .A1(n3340), .A2(n3459), .B1(\RegFilePlugin_regFile[19][14] ), .B2(n3340), .Z(n4826) );
  aoim22d1 U5458 ( .A1(n3347), .A2(n3485), .B1(\RegFilePlugin_regFile[19][13] ), .B2(n3346), .Z(n4825) );
  aoim22d1 U5459 ( .A1(n3346), .A2(n3460), .B1(\RegFilePlugin_regFile[19][12] ), .B2(n3340), .Z(n4824) );
  aoim22d1 U5460 ( .A1(n3347), .A2(n3461), .B1(\RegFilePlugin_regFile[19][11] ), .B2(n3345), .Z(n4823) );
  aoim22d1 U5461 ( .A1(n3347), .A2(n3462), .B1(\RegFilePlugin_regFile[19][10] ), .B2(n3345), .Z(n4822) );
  aoim22d1 U5462 ( .A1(n3345), .A2(n3463), .B1(\RegFilePlugin_regFile[19][9] ), 
        .B2(n3345), .Z(n4821) );
  aoim22d1 U5463 ( .A1(n3347), .A2(n3541), .B1(\RegFilePlugin_regFile[19][8] ), 
        .B2(n3345), .Z(n4820) );
  aoim22d1 U5464 ( .A1(n3340), .A2(n3543), .B1(\RegFilePlugin_regFile[19][7] ), 
        .B2(n3345), .Z(n4819) );
  aoim22d1 U5465 ( .A1(n3347), .A2(n3467), .B1(\RegFilePlugin_regFile[19][6] ), 
        .B2(n3345), .Z(n4818) );
  aoim22d1 U5466 ( .A1(n3347), .A2(n3468), .B1(\RegFilePlugin_regFile[19][5] ), 
        .B2(n3347), .Z(n4817) );
  aoim22d1 U5467 ( .A1(n3346), .A2(n3469), .B1(\RegFilePlugin_regFile[19][4] ), 
        .B2(n3347), .Z(n4816) );
  aoim22d1 U5468 ( .A1(n3340), .A2(n3551), .B1(\RegFilePlugin_regFile[19][3] ), 
        .B2(n3347), .Z(n4815) );
  aoim22d1 U5469 ( .A1(n3347), .A2(n3472), .B1(\RegFilePlugin_regFile[19][2] ), 
        .B2(n3347), .Z(n4814) );
  aoim22d1 U5470 ( .A1(n3347), .A2(n3554), .B1(\RegFilePlugin_regFile[19][1] ), 
        .B2(n3347), .Z(n4813) );
  nr02d1 U5471 ( .A1(n3481), .A2(n3356), .ZN(n3348) );
  buffd1 U5472 ( .I(n3348), .Z(n3350) );
  aoim22d1 U5473 ( .A1(n3350), .A2(n3500), .B1(\RegFilePlugin_regFile[18][0] ), 
        .B2(n3348), .Z(n4812) );
  buffd1 U5474 ( .I(n3348), .Z(n3349) );
  aoim22d1 U5475 ( .A1(n3349), .A2(n3338), .B1(\RegFilePlugin_regFile[18][31] ), .B2(n3351), .Z(n4811) );
  aoim22d1 U5476 ( .A1(n3350), .A2(n3503), .B1(\RegFilePlugin_regFile[18][30] ), .B2(n3349), .Z(n4810) );
  aoim22d1 U5477 ( .A1(n3350), .A2(n3505), .B1(\RegFilePlugin_regFile[18][29] ), .B2(n3349), .Z(n4809) );
  buffd1 U5478 ( .I(n3348), .Z(n3351) );
  aoim22d1 U5479 ( .A1(n3351), .A2(n3484), .B1(\RegFilePlugin_regFile[18][28] ), .B2(n3349), .Z(n4808) );
  aoim22d1 U5480 ( .A1(n3350), .A2(n3508), .B1(\RegFilePlugin_regFile[18][27] ), .B2(n3351), .Z(n4807) );
  aoim22d1 U5481 ( .A1(n3350), .A2(n3510), .B1(\RegFilePlugin_regFile[18][26] ), .B2(n3349), .Z(n4806) );
  aoim22d1 U5482 ( .A1(n3349), .A2(n3512), .B1(\RegFilePlugin_regFile[18][25] ), .B2(n3351), .Z(n4805) );
  aoim22d1 U5483 ( .A1(n3349), .A2(n3341), .B1(\RegFilePlugin_regFile[18][24] ), .B2(n3350), .Z(n4804) );
  aoim22d1 U5484 ( .A1(n3350), .A2(n3454), .B1(\RegFilePlugin_regFile[18][23] ), .B2(n3351), .Z(n4803) );
  aoim22d1 U5485 ( .A1(n3350), .A2(n3517), .B1(\RegFilePlugin_regFile[18][22] ), .B2(n3350), .Z(n4802) );
  aoim22d1 U5486 ( .A1(n3350), .A2(n3519), .B1(\RegFilePlugin_regFile[18][21] ), .B2(n3350), .Z(n4801) );
  aoim22d1 U5487 ( .A1(n3349), .A2(n3521), .B1(\RegFilePlugin_regFile[18][20] ), .B2(n3351), .Z(n4800) );
  aoim22d1 U5488 ( .A1(n3351), .A2(n3344), .B1(\RegFilePlugin_regFile[18][19] ), .B2(n3350), .Z(n4799) );
  aoim22d1 U5489 ( .A1(n3348), .A2(n3456), .B1(\RegFilePlugin_regFile[18][18] ), .B2(n3350), .Z(n4798) );
  aoim22d1 U5490 ( .A1(n3351), .A2(n3527), .B1(\RegFilePlugin_regFile[18][17] ), .B2(n3351), .Z(n4797) );
  aoim22d1 U5491 ( .A1(n3350), .A2(n3458), .B1(\RegFilePlugin_regFile[18][16] ), .B2(n3351), .Z(n4796) );
  aoim22d1 U5492 ( .A1(n3349), .A2(n3366), .B1(\RegFilePlugin_regFile[18][15] ), .B2(n3351), .Z(n4795) );
  aoim22d1 U5493 ( .A1(n3351), .A2(n3459), .B1(\RegFilePlugin_regFile[18][14] ), .B2(n3351), .Z(n4794) );
  aoim22d1 U5494 ( .A1(n3348), .A2(n3485), .B1(\RegFilePlugin_regFile[18][13] ), .B2(n3351), .Z(n4793) );
  aoim22d1 U5495 ( .A1(n3350), .A2(n3460), .B1(\RegFilePlugin_regFile[18][12] ), .B2(n3351), .Z(n4792) );
  aoim22d1 U5496 ( .A1(n3349), .A2(n3461), .B1(\RegFilePlugin_regFile[18][11] ), .B2(n3349), .Z(n4791) );
  aoim22d1 U5497 ( .A1(n3348), .A2(n3462), .B1(\RegFilePlugin_regFile[18][10] ), .B2(n3349), .Z(n4790) );
  aoim22d1 U5498 ( .A1(n3349), .A2(n3463), .B1(\RegFilePlugin_regFile[18][9] ), 
        .B2(n3349), .Z(n4789) );
  aoim22d1 U5499 ( .A1(n3348), .A2(n3464), .B1(\RegFilePlugin_regFile[18][8] ), 
        .B2(n3349), .Z(n4788) );
  aoim22d1 U5500 ( .A1(n3351), .A2(n3465), .B1(\RegFilePlugin_regFile[18][7] ), 
        .B2(n3349), .Z(n4787) );
  aoim22d1 U5501 ( .A1(n3348), .A2(n3467), .B1(\RegFilePlugin_regFile[18][6] ), 
        .B2(n3349), .Z(n4786) );
  aoim22d1 U5502 ( .A1(n3348), .A2(n3468), .B1(\RegFilePlugin_regFile[18][5] ), 
        .B2(n3348), .Z(n4785) );
  aoim22d1 U5503 ( .A1(n3350), .A2(n3469), .B1(\RegFilePlugin_regFile[18][4] ), 
        .B2(n3350), .Z(n4784) );
  aoim22d1 U5504 ( .A1(n3351), .A2(n3471), .B1(\RegFilePlugin_regFile[18][3] ), 
        .B2(n3348), .Z(n4783) );
  aoim22d1 U5505 ( .A1(n3348), .A2(n3472), .B1(\RegFilePlugin_regFile[18][2] ), 
        .B2(n3348), .Z(n4782) );
  aoim22d1 U5506 ( .A1(n3348), .A2(n3473), .B1(\RegFilePlugin_regFile[18][1] ), 
        .B2(n3348), .Z(n4781) );
  nr02d1 U5507 ( .A1(n3489), .A2(n3356), .ZN(n3352) );
  buffd1 U5508 ( .I(n3352), .Z(n3354) );
  buffd1 U5509 ( .I(n3352), .Z(n3355) );
  aoim22d1 U5510 ( .A1(n3354), .A2(n3500), .B1(\RegFilePlugin_regFile[17][0] ), 
        .B2(n3355), .Z(n4780) );
  buffd1 U5511 ( .I(n3352), .Z(n3353) );
  aoim22d1 U5512 ( .A1(n3353), .A2(n3450), .B1(\RegFilePlugin_regFile[17][31] ), .B2(n3355), .Z(n4779) );
  aoim22d1 U5513 ( .A1(n3354), .A2(n3503), .B1(\RegFilePlugin_regFile[17][30] ), .B2(n3353), .Z(n4778) );
  aoim22d1 U5514 ( .A1(n3354), .A2(n3339), .B1(\RegFilePlugin_regFile[17][29] ), .B2(n3353), .Z(n4777) );
  aoim22d1 U5515 ( .A1(n3352), .A2(n3484), .B1(\RegFilePlugin_regFile[17][28] ), .B2(n3353), .Z(n4776) );
  aoim22d1 U5516 ( .A1(n3354), .A2(n3508), .B1(\RegFilePlugin_regFile[17][27] ), .B2(n3352), .Z(n4775) );
  aoim22d1 U5517 ( .A1(n3354), .A2(n3510), .B1(\RegFilePlugin_regFile[17][26] ), .B2(n3353), .Z(n4774) );
  aoim22d1 U5518 ( .A1(n3353), .A2(n3512), .B1(\RegFilePlugin_regFile[17][25] ), .B2(n3354), .Z(n4773) );
  aoim22d1 U5519 ( .A1(n3353), .A2(n3453), .B1(\RegFilePlugin_regFile[17][24] ), .B2(n3354), .Z(n4772) );
  aoim22d1 U5520 ( .A1(n3354), .A2(n3454), .B1(\RegFilePlugin_regFile[17][23] ), .B2(n3352), .Z(n4771) );
  aoim22d1 U5521 ( .A1(n3354), .A2(n3517), .B1(\RegFilePlugin_regFile[17][22] ), .B2(n3354), .Z(n4770) );
  aoim22d1 U5522 ( .A1(n3354), .A2(n3342), .B1(\RegFilePlugin_regFile[17][21] ), .B2(n3354), .Z(n4769) );
  aoim22d1 U5523 ( .A1(n3353), .A2(n3343), .B1(\RegFilePlugin_regFile[17][20] ), .B2(n3352), .Z(n4768) );
  aoim22d1 U5524 ( .A1(n3352), .A2(n3523), .B1(\RegFilePlugin_regFile[17][19] ), .B2(n3354), .Z(n4767) );
  aoim22d1 U5525 ( .A1(n3355), .A2(n3456), .B1(\RegFilePlugin_regFile[17][18] ), .B2(n3354), .Z(n4766) );
  aoim22d1 U5526 ( .A1(n3355), .A2(n3527), .B1(\RegFilePlugin_regFile[17][17] ), .B2(n3353), .Z(n4765) );
  aoim22d1 U5527 ( .A1(n3354), .A2(n3529), .B1(\RegFilePlugin_regFile[17][16] ), .B2(n3352), .Z(n4764) );
  aoim22d1 U5528 ( .A1(n3353), .A2(n3366), .B1(\RegFilePlugin_regFile[17][15] ), .B2(n3352), .Z(n4763) );
  aoim22d1 U5529 ( .A1(n3352), .A2(n3459), .B1(\RegFilePlugin_regFile[17][14] ), .B2(n3352), .Z(n4762) );
  aoim22d1 U5530 ( .A1(n3355), .A2(n3485), .B1(\RegFilePlugin_regFile[17][13] ), .B2(n3352), .Z(n4761) );
  aoim22d1 U5531 ( .A1(n3354), .A2(n3460), .B1(\RegFilePlugin_regFile[17][12] ), .B2(n3352), .Z(n4760) );
  aoim22d1 U5532 ( .A1(n3355), .A2(n3461), .B1(\RegFilePlugin_regFile[17][11] ), .B2(n3353), .Z(n4759) );
  aoim22d1 U5533 ( .A1(n3355), .A2(n3462), .B1(\RegFilePlugin_regFile[17][10] ), .B2(n3353), .Z(n4758) );
  aoim22d1 U5534 ( .A1(n3353), .A2(n3463), .B1(\RegFilePlugin_regFile[17][9] ), 
        .B2(n3353), .Z(n4757) );
  aoim22d1 U5535 ( .A1(n3355), .A2(n3541), .B1(\RegFilePlugin_regFile[17][8] ), 
        .B2(n3353), .Z(n4756) );
  aoim22d1 U5536 ( .A1(n3352), .A2(n3543), .B1(\RegFilePlugin_regFile[17][7] ), 
        .B2(n3353), .Z(n4755) );
  aoim22d1 U5537 ( .A1(n3355), .A2(n3467), .B1(\RegFilePlugin_regFile[17][6] ), 
        .B2(n3353), .Z(n4754) );
  aoim22d1 U5538 ( .A1(n3355), .A2(n3468), .B1(\RegFilePlugin_regFile[17][5] ), 
        .B2(n3355), .Z(n4753) );
  aoim22d1 U5539 ( .A1(n3354), .A2(n3469), .B1(\RegFilePlugin_regFile[17][4] ), 
        .B2(n3355), .Z(n4752) );
  aoim22d1 U5540 ( .A1(n3352), .A2(n3551), .B1(\RegFilePlugin_regFile[17][3] ), 
        .B2(n3355), .Z(n4751) );
  aoim22d1 U5541 ( .A1(n3355), .A2(n3472), .B1(\RegFilePlugin_regFile[17][2] ), 
        .B2(n3355), .Z(n4750) );
  aoim22d1 U5542 ( .A1(n3355), .A2(n3554), .B1(\RegFilePlugin_regFile[17][1] ), 
        .B2(n3355), .Z(n4749) );
  nr02d1 U5543 ( .A1(n3498), .A2(n3356), .ZN(n3357) );
  buffd1 U5544 ( .I(n3357), .Z(n3359) );
  buffd1 U5545 ( .I(n3357), .Z(n3360) );
  aoim22d1 U5546 ( .A1(n3359), .A2(n3500), .B1(\RegFilePlugin_regFile[16][0] ), 
        .B2(n3360), .Z(n4748) );
  buffd1 U5547 ( .I(n3357), .Z(n3358) );
  aoim22d1 U5548 ( .A1(n3358), .A2(n3338), .B1(\RegFilePlugin_regFile[16][31] ), .B2(n3360), .Z(n4747) );
  aoim22d1 U5549 ( .A1(n3359), .A2(n3503), .B1(\RegFilePlugin_regFile[16][30] ), .B2(n3358), .Z(n4746) );
  aoim22d1 U5550 ( .A1(n3359), .A2(n3505), .B1(\RegFilePlugin_regFile[16][29] ), .B2(n3358), .Z(n4745) );
  aoim22d1 U5551 ( .A1(n3357), .A2(n3484), .B1(\RegFilePlugin_regFile[16][28] ), .B2(n3358), .Z(n4744) );
  aoim22d1 U5552 ( .A1(n3359), .A2(n3508), .B1(\RegFilePlugin_regFile[16][27] ), .B2(n3357), .Z(n4743) );
  aoim22d1 U5553 ( .A1(n3359), .A2(n3510), .B1(\RegFilePlugin_regFile[16][26] ), .B2(n3358), .Z(n4742) );
  aoim22d1 U5554 ( .A1(n3358), .A2(n3512), .B1(\RegFilePlugin_regFile[16][25] ), .B2(n3357), .Z(n4741) );
  aoim22d1 U5555 ( .A1(n3358), .A2(n3341), .B1(\RegFilePlugin_regFile[16][24] ), .B2(n3359), .Z(n4740) );
  aoim22d1 U5556 ( .A1(n3359), .A2(n3454), .B1(\RegFilePlugin_regFile[16][23] ), .B2(n3357), .Z(n4739) );
  aoim22d1 U5557 ( .A1(n3359), .A2(n3517), .B1(\RegFilePlugin_regFile[16][22] ), .B2(n3359), .Z(n4738) );
  aoim22d1 U5558 ( .A1(n3359), .A2(n3519), .B1(\RegFilePlugin_regFile[16][21] ), .B2(n3359), .Z(n4737) );
  aoim22d1 U5559 ( .A1(n3358), .A2(n3521), .B1(\RegFilePlugin_regFile[16][20] ), .B2(n3357), .Z(n4736) );
  aoim22d1 U5560 ( .A1(n3357), .A2(n3523), .B1(\RegFilePlugin_regFile[16][19] ), .B2(n3359), .Z(n4735) );
  aoim22d1 U5561 ( .A1(n3360), .A2(n3456), .B1(\RegFilePlugin_regFile[16][18] ), .B2(n3359), .Z(n4734) );
  aoim22d1 U5562 ( .A1(n3360), .A2(n3527), .B1(\RegFilePlugin_regFile[16][17] ), .B2(n3359), .Z(n4733) );
  aoim22d1 U5563 ( .A1(n3359), .A2(n3458), .B1(\RegFilePlugin_regFile[16][16] ), .B2(n3358), .Z(n4732) );
  aoim22d1 U5564 ( .A1(n3358), .A2(n3366), .B1(\RegFilePlugin_regFile[16][15] ), .B2(n3357), .Z(n4731) );
  aoim22d1 U5565 ( .A1(n3357), .A2(n3459), .B1(\RegFilePlugin_regFile[16][14] ), .B2(n3357), .Z(n4730) );
  aoim22d1 U5566 ( .A1(n3360), .A2(n3485), .B1(\RegFilePlugin_regFile[16][13] ), .B2(n3357), .Z(n4729) );
  aoim22d1 U5567 ( .A1(n3359), .A2(n3460), .B1(\RegFilePlugin_regFile[16][12] ), .B2(n3357), .Z(n4728) );
  aoim22d1 U5568 ( .A1(n3360), .A2(n3461), .B1(\RegFilePlugin_regFile[16][11] ), .B2(n3358), .Z(n4727) );
  aoim22d1 U5569 ( .A1(n3360), .A2(n3462), .B1(\RegFilePlugin_regFile[16][10] ), .B2(n3358), .Z(n4726) );
  aoim22d1 U5570 ( .A1(n3358), .A2(n3463), .B1(\RegFilePlugin_regFile[16][9] ), 
        .B2(n3358), .Z(n4725) );
  aoim22d1 U5571 ( .A1(n3360), .A2(n3464), .B1(\RegFilePlugin_regFile[16][8] ), 
        .B2(n3358), .Z(n4724) );
  aoim22d1 U5572 ( .A1(n3357), .A2(n3465), .B1(\RegFilePlugin_regFile[16][7] ), 
        .B2(n3358), .Z(n4723) );
  aoim22d1 U5573 ( .A1(n3360), .A2(n3467), .B1(\RegFilePlugin_regFile[16][6] ), 
        .B2(n3358), .Z(n4722) );
  aoim22d1 U5574 ( .A1(n3360), .A2(n3468), .B1(\RegFilePlugin_regFile[16][5] ), 
        .B2(n3360), .Z(n4721) );
  aoim22d1 U5575 ( .A1(n3359), .A2(n3469), .B1(\RegFilePlugin_regFile[16][4] ), 
        .B2(n3360), .Z(n4720) );
  aoim22d1 U5576 ( .A1(n3357), .A2(n3471), .B1(\RegFilePlugin_regFile[16][3] ), 
        .B2(n3360), .Z(n4719) );
  aoim22d1 U5577 ( .A1(n3360), .A2(n3472), .B1(\RegFilePlugin_regFile[16][2] ), 
        .B2(n3360), .Z(n4718) );
  aoim22d1 U5578 ( .A1(n3360), .A2(n3473), .B1(\RegFilePlugin_regFile[16][1] ), 
        .B2(n3360), .Z(n4717) );
  inv0d0 U5579 ( .I(_zz_lastStageRegFileWrite_payload_address[11]), .ZN(n3431)
         );
  nd03d0 U5580 ( .A1(_zz_lastStageRegFileWrite_payload_address[10]), .A2(n3433), .A3(n3431), .ZN(n3392) );
  nr02d1 U5581 ( .A1(n3434), .A2(n3392), .ZN(n3361) );
  buffd1 U5582 ( .I(n3361), .Z(n3364) );
  aoim22d1 U5583 ( .A1(n3361), .A2(n3500), .B1(\RegFilePlugin_regFile[15][0] ), 
        .B2(n3364), .Z(n4716) );
  buffd1 U5584 ( .I(n3361), .Z(n3362) );
  aoim22d1 U5585 ( .A1(n3362), .A2(n3338), .B1(\RegFilePlugin_regFile[15][31] ), .B2(n3364), .Z(n4715) );
  aoim22d1 U5586 ( .A1(n3363), .A2(n3503), .B1(\RegFilePlugin_regFile[15][30] ), .B2(n3362), .Z(n4714) );
  aoim22d1 U5587 ( .A1(n3361), .A2(n3505), .B1(\RegFilePlugin_regFile[15][29] ), .B2(n3362), .Z(n4713) );
  buffd1 U5588 ( .I(n3361), .Z(n3363) );
  aoim22d1 U5589 ( .A1(n3363), .A2(n3484), .B1(\RegFilePlugin_regFile[15][28] ), .B2(n3362), .Z(n4712) );
  aoim22d1 U5590 ( .A1(n3361), .A2(n3508), .B1(\RegFilePlugin_regFile[15][27] ), .B2(n3363), .Z(n4711) );
  aoim22d1 U5591 ( .A1(n3361), .A2(n3510), .B1(\RegFilePlugin_regFile[15][26] ), .B2(n3362), .Z(n4710) );
  aoim22d1 U5592 ( .A1(n3362), .A2(n3512), .B1(\RegFilePlugin_regFile[15][25] ), .B2(n3363), .Z(n4709) );
  aoim22d1 U5593 ( .A1(n3362), .A2(n3341), .B1(\RegFilePlugin_regFile[15][24] ), .B2(n3361), .Z(n4708) );
  aoim22d1 U5594 ( .A1(n3364), .A2(n3454), .B1(\RegFilePlugin_regFile[15][23] ), .B2(n3363), .Z(n4707) );
  aoim22d1 U5595 ( .A1(n3361), .A2(n3517), .B1(\RegFilePlugin_regFile[15][22] ), .B2(n3361), .Z(n4706) );
  aoim22d1 U5596 ( .A1(n3361), .A2(n3519), .B1(\RegFilePlugin_regFile[15][21] ), .B2(n3361), .Z(n4705) );
  aoim22d1 U5597 ( .A1(n3362), .A2(n3521), .B1(\RegFilePlugin_regFile[15][20] ), .B2(n3363), .Z(n4704) );
  aoim22d1 U5598 ( .A1(n3363), .A2(n3523), .B1(\RegFilePlugin_regFile[15][19] ), .B2(n3361), .Z(n4703) );
  aoim22d1 U5599 ( .A1(n3364), .A2(n3456), .B1(\RegFilePlugin_regFile[15][18] ), .B2(n3361), .Z(n4702) );
  aoim22d1 U5600 ( .A1(n3363), .A2(n3527), .B1(\RegFilePlugin_regFile[15][17] ), .B2(n3363), .Z(n4701) );
  aoim22d1 U5601 ( .A1(n3362), .A2(n3529), .B1(\RegFilePlugin_regFile[15][16] ), .B2(n3363), .Z(n4700) );
  aoim22d1 U5602 ( .A1(n3362), .A2(n3366), .B1(\RegFilePlugin_regFile[15][15] ), .B2(n3363), .Z(n4699) );
  aoim22d1 U5603 ( .A1(n3363), .A2(n3459), .B1(\RegFilePlugin_regFile[15][14] ), .B2(n3363), .Z(n4698) );
  aoim22d1 U5604 ( .A1(n3364), .A2(n3534), .B1(\RegFilePlugin_regFile[15][13] ), .B2(n3363), .Z(n4697) );
  aoim22d1 U5605 ( .A1(n3361), .A2(n3460), .B1(\RegFilePlugin_regFile[15][12] ), .B2(n3363), .Z(n4696) );
  aoim22d1 U5606 ( .A1(n3364), .A2(n3461), .B1(\RegFilePlugin_regFile[15][11] ), .B2(n3362), .Z(n4695) );
  aoim22d1 U5607 ( .A1(n3364), .A2(n3462), .B1(\RegFilePlugin_regFile[15][10] ), .B2(n3362), .Z(n4694) );
  aoim22d1 U5608 ( .A1(n3362), .A2(n3463), .B1(\RegFilePlugin_regFile[15][9] ), 
        .B2(n3362), .Z(n4693) );
  aoim22d1 U5609 ( .A1(n3364), .A2(n3541), .B1(\RegFilePlugin_regFile[15][8] ), 
        .B2(n3362), .Z(n4692) );
  aoim22d1 U5610 ( .A1(n3363), .A2(n3543), .B1(\RegFilePlugin_regFile[15][7] ), 
        .B2(n3362), .Z(n4691) );
  aoim22d1 U5611 ( .A1(n3364), .A2(n3467), .B1(\RegFilePlugin_regFile[15][6] ), 
        .B2(n3362), .Z(n4690) );
  aoim22d1 U5612 ( .A1(n3364), .A2(n3468), .B1(\RegFilePlugin_regFile[15][5] ), 
        .B2(n3364), .Z(n4689) );
  aoim22d1 U5613 ( .A1(n3361), .A2(n3469), .B1(\RegFilePlugin_regFile[15][4] ), 
        .B2(n3364), .Z(n4688) );
  aoim22d1 U5614 ( .A1(n3363), .A2(n3551), .B1(\RegFilePlugin_regFile[15][3] ), 
        .B2(n3364), .Z(n4687) );
  aoim22d1 U5615 ( .A1(n3364), .A2(n3472), .B1(\RegFilePlugin_regFile[15][2] ), 
        .B2(n3364), .Z(n4686) );
  aoim22d1 U5616 ( .A1(n3364), .A2(n3554), .B1(\RegFilePlugin_regFile[15][1] ), 
        .B2(n3364), .Z(n4685) );
  nr02d1 U5617 ( .A1(n3439), .A2(n3392), .ZN(n3365) );
  buffd1 U5618 ( .I(n3365), .Z(n3368) );
  buffd1 U5619 ( .I(n3365), .Z(n3369) );
  aoim22d1 U5620 ( .A1(n3368), .A2(n3500), .B1(\RegFilePlugin_regFile[14][0] ), 
        .B2(n3369), .Z(n4684) );
  buffd1 U5621 ( .I(n3365), .Z(n3367) );
  aoim22d1 U5622 ( .A1(n3367), .A2(n3338), .B1(\RegFilePlugin_regFile[14][31] ), .B2(n3369), .Z(n4683) );
  aoim22d1 U5623 ( .A1(n3368), .A2(n3503), .B1(\RegFilePlugin_regFile[14][30] ), .B2(n3367), .Z(n4682) );
  aoim22d1 U5624 ( .A1(n3368), .A2(n3505), .B1(\RegFilePlugin_regFile[14][29] ), .B2(n3367), .Z(n4681) );
  aoim22d1 U5625 ( .A1(n3365), .A2(n3484), .B1(\RegFilePlugin_regFile[14][28] ), .B2(n3367), .Z(n4680) );
  aoim22d1 U5626 ( .A1(n3368), .A2(n3508), .B1(\RegFilePlugin_regFile[14][27] ), .B2(n3365), .Z(n4679) );
  aoim22d1 U5627 ( .A1(n3368), .A2(n3510), .B1(\RegFilePlugin_regFile[14][26] ), .B2(n3367), .Z(n4678) );
  aoim22d1 U5628 ( .A1(n3367), .A2(n3512), .B1(\RegFilePlugin_regFile[14][25] ), .B2(n3365), .Z(n4677) );
  aoim22d1 U5629 ( .A1(n3367), .A2(n3341), .B1(\RegFilePlugin_regFile[14][24] ), .B2(n3368), .Z(n4676) );
  aoim22d1 U5630 ( .A1(n3368), .A2(n3454), .B1(\RegFilePlugin_regFile[14][23] ), .B2(n3365), .Z(n4675) );
  aoim22d1 U5631 ( .A1(n3368), .A2(n3517), .B1(\RegFilePlugin_regFile[14][22] ), .B2(n3368), .Z(n4674) );
  aoim22d1 U5632 ( .A1(n3368), .A2(n3519), .B1(\RegFilePlugin_regFile[14][21] ), .B2(n3368), .Z(n4673) );
  aoim22d1 U5633 ( .A1(n3367), .A2(n3521), .B1(\RegFilePlugin_regFile[14][20] ), .B2(n3365), .Z(n4672) );
  aoim22d1 U5634 ( .A1(n3365), .A2(n3523), .B1(\RegFilePlugin_regFile[14][19] ), .B2(n3368), .Z(n4671) );
  aoim22d1 U5635 ( .A1(n3369), .A2(n3456), .B1(\RegFilePlugin_regFile[14][18] ), .B2(n3368), .Z(n4670) );
  aoim22d1 U5636 ( .A1(n3365), .A2(n3527), .B1(\RegFilePlugin_regFile[14][17] ), .B2(n3368), .Z(n4669) );
  aoim22d1 U5637 ( .A1(n3368), .A2(n3529), .B1(\RegFilePlugin_regFile[14][16] ), .B2(n3367), .Z(n4668) );
  aoim22d1 U5638 ( .A1(n3367), .A2(n3366), .B1(\RegFilePlugin_regFile[14][15] ), .B2(n3365), .Z(n4667) );
  aoim22d1 U5639 ( .A1(n3365), .A2(n3459), .B1(\RegFilePlugin_regFile[14][14] ), .B2(n3365), .Z(n4666) );
  aoim22d1 U5640 ( .A1(n3369), .A2(n3534), .B1(\RegFilePlugin_regFile[14][13] ), .B2(n3369), .Z(n4665) );
  aoim22d1 U5641 ( .A1(n3368), .A2(n3460), .B1(\RegFilePlugin_regFile[14][12] ), .B2(n3365), .Z(n4664) );
  aoim22d1 U5642 ( .A1(n3369), .A2(n3461), .B1(\RegFilePlugin_regFile[14][11] ), .B2(n3367), .Z(n4663) );
  aoim22d1 U5643 ( .A1(n3369), .A2(n3462), .B1(\RegFilePlugin_regFile[14][10] ), .B2(n3367), .Z(n4662) );
  aoim22d1 U5644 ( .A1(n3367), .A2(n3463), .B1(\RegFilePlugin_regFile[14][9] ), 
        .B2(n3367), .Z(n4661) );
  aoim22d1 U5645 ( .A1(n3369), .A2(n3541), .B1(\RegFilePlugin_regFile[14][8] ), 
        .B2(n3367), .Z(n4660) );
  aoim22d1 U5646 ( .A1(n3365), .A2(n3543), .B1(\RegFilePlugin_regFile[14][7] ), 
        .B2(n3367), .Z(n4659) );
  aoim22d1 U5647 ( .A1(n3369), .A2(n3467), .B1(\RegFilePlugin_regFile[14][6] ), 
        .B2(n3367), .Z(n4658) );
  aoim22d1 U5648 ( .A1(n3369), .A2(n3468), .B1(\RegFilePlugin_regFile[14][5] ), 
        .B2(n3369), .Z(n4657) );
  aoim22d1 U5649 ( .A1(n3368), .A2(n3469), .B1(\RegFilePlugin_regFile[14][4] ), 
        .B2(n3369), .Z(n4656) );
  aoim22d1 U5650 ( .A1(n3365), .A2(n3551), .B1(\RegFilePlugin_regFile[14][3] ), 
        .B2(n3369), .Z(n4655) );
  aoim22d1 U5651 ( .A1(n3369), .A2(n3472), .B1(\RegFilePlugin_regFile[14][2] ), 
        .B2(n3369), .Z(n4654) );
  aoim22d1 U5652 ( .A1(n3369), .A2(n3554), .B1(\RegFilePlugin_regFile[14][1] ), 
        .B2(n3369), .Z(n4653) );
  buffd1 U5653 ( .I(n3370), .Z(n3372) );
  buffd1 U5654 ( .I(n3370), .Z(n3374) );
  aoim22d1 U5655 ( .A1(n3372), .A2(n3482), .B1(\RegFilePlugin_regFile[13][0] ), 
        .B2(n3374), .Z(n4652) );
  buffd1 U5656 ( .I(n3370), .Z(n3371) );
  aoim22d1 U5657 ( .A1(n3371), .A2(n3450), .B1(\RegFilePlugin_regFile[13][31] ), .B2(n3374), .Z(n4651) );
  aoim22d1 U5658 ( .A1(n3372), .A2(n3490), .B1(\RegFilePlugin_regFile[13][30] ), .B2(n3371), .Z(n4650) );
  aoim22d1 U5659 ( .A1(n3372), .A2(n3339), .B1(\RegFilePlugin_regFile[13][29] ), .B2(n3371), .Z(n4649) );
  buffd1 U5660 ( .I(n3370), .Z(n3373) );
  aoim22d1 U5661 ( .A1(n3373), .A2(n3476), .B1(\RegFilePlugin_regFile[13][28] ), .B2(n3371), .Z(n4648) );
  aoim22d1 U5662 ( .A1(n3372), .A2(n3492), .B1(\RegFilePlugin_regFile[13][27] ), .B2(n3373), .Z(n4647) );
  aoim22d1 U5663 ( .A1(n3372), .A2(n3493), .B1(\RegFilePlugin_regFile[13][26] ), .B2(n3371), .Z(n4646) );
  aoim22d1 U5664 ( .A1(n3371), .A2(n3452), .B1(\RegFilePlugin_regFile[13][25] ), .B2(n3373), .Z(n4645) );
  aoim22d1 U5665 ( .A1(n3371), .A2(n3453), .B1(\RegFilePlugin_regFile[13][24] ), .B2(n3372), .Z(n4644) );
  aoim22d1 U5666 ( .A1(n3372), .A2(n3454), .B1(\RegFilePlugin_regFile[13][23] ), .B2(n3373), .Z(n4643) );
  aoim22d1 U5667 ( .A1(n3372), .A2(n3455), .B1(\RegFilePlugin_regFile[13][22] ), .B2(n3372), .Z(n4642) );
  aoim22d1 U5668 ( .A1(n3372), .A2(n3342), .B1(\RegFilePlugin_regFile[13][21] ), .B2(n3372), .Z(n4641) );
  aoim22d1 U5669 ( .A1(n3371), .A2(n3343), .B1(\RegFilePlugin_regFile[13][20] ), .B2(n3373), .Z(n4640) );
  aoim22d1 U5670 ( .A1(n3373), .A2(n3344), .B1(\RegFilePlugin_regFile[13][19] ), .B2(n3372), .Z(n4639) );
  aoim22d1 U5671 ( .A1(n3374), .A2(n3456), .B1(\RegFilePlugin_regFile[13][18] ), .B2(n3372), .Z(n4638) );
  aoim22d1 U5672 ( .A1(n3373), .A2(n3457), .B1(\RegFilePlugin_regFile[13][17] ), .B2(n3373), .Z(n4637) );
  aoim22d1 U5673 ( .A1(n3372), .A2(n3458), .B1(\RegFilePlugin_regFile[13][16] ), .B2(n3373), .Z(n4636) );
  aoim22d1 U5674 ( .A1(n3371), .A2(n3531), .B1(\RegFilePlugin_regFile[13][15] ), .B2(n3373), .Z(n4635) );
  aoim22d1 U5675 ( .A1(n3373), .A2(n3459), .B1(\RegFilePlugin_regFile[13][14] ), .B2(n3373), .Z(n4634) );
  aoim22d1 U5676 ( .A1(n3374), .A2(n3534), .B1(\RegFilePlugin_regFile[13][13] ), .B2(n3373), .Z(n4633) );
  aoim22d1 U5677 ( .A1(n3372), .A2(n3460), .B1(\RegFilePlugin_regFile[13][12] ), .B2(n3373), .Z(n4632) );
  aoim22d1 U5678 ( .A1(n3374), .A2(n3461), .B1(\RegFilePlugin_regFile[13][11] ), .B2(n3371), .Z(n4631) );
  aoim22d1 U5679 ( .A1(n3374), .A2(n3462), .B1(\RegFilePlugin_regFile[13][10] ), .B2(n3371), .Z(n4630) );
  aoim22d1 U5680 ( .A1(n3371), .A2(n3463), .B1(\RegFilePlugin_regFile[13][9] ), 
        .B2(n3371), .Z(n4629) );
  aoim22d1 U5681 ( .A1(n3374), .A2(n3464), .B1(\RegFilePlugin_regFile[13][8] ), 
        .B2(n3371), .Z(n4628) );
  aoim22d1 U5682 ( .A1(n3373), .A2(n3465), .B1(\RegFilePlugin_regFile[13][7] ), 
        .B2(n3371), .Z(n4627) );
  aoim22d1 U5683 ( .A1(n3374), .A2(n3467), .B1(\RegFilePlugin_regFile[13][6] ), 
        .B2(n3371), .Z(n4626) );
  aoim22d1 U5684 ( .A1(n3374), .A2(n3468), .B1(\RegFilePlugin_regFile[13][5] ), 
        .B2(n3374), .Z(n4625) );
  aoim22d1 U5685 ( .A1(n3372), .A2(n3469), .B1(\RegFilePlugin_regFile[13][4] ), 
        .B2(n3374), .Z(n4624) );
  aoim22d1 U5686 ( .A1(n3373), .A2(n3471), .B1(\RegFilePlugin_regFile[13][3] ), 
        .B2(n3374), .Z(n4623) );
  aoim22d1 U5687 ( .A1(n3374), .A2(n3472), .B1(\RegFilePlugin_regFile[13][2] ), 
        .B2(n3374), .Z(n4622) );
  aoim22d1 U5688 ( .A1(n3374), .A2(n3473), .B1(\RegFilePlugin_regFile[13][1] ), 
        .B2(n3374), .Z(n4621) );
  nr02d1 U5689 ( .A1(n3449), .A2(n3392), .ZN(n3375) );
  buffd1 U5690 ( .I(n3375), .Z(n3376) );
  buffd1 U5691 ( .I(n3375), .Z(n3378) );
  aoim22d1 U5692 ( .A1(n3376), .A2(n3482), .B1(\RegFilePlugin_regFile[12][0] ), 
        .B2(n3378), .Z(n4620) );
  aoim22d1 U5693 ( .A1(n3377), .A2(n3450), .B1(\RegFilePlugin_regFile[12][31] ), .B2(n3378), .Z(n4619) );
  aoim22d1 U5694 ( .A1(n3376), .A2(n3490), .B1(\RegFilePlugin_regFile[12][30] ), .B2(n3375), .Z(n4618) );
  aoim22d1 U5695 ( .A1(n3376), .A2(n3339), .B1(\RegFilePlugin_regFile[12][29] ), .B2(n3375), .Z(n4617) );
  buffd1 U5696 ( .I(n3375), .Z(n3377) );
  aoim22d1 U5697 ( .A1(n3377), .A2(n3476), .B1(\RegFilePlugin_regFile[12][28] ), .B2(n3375), .Z(n4616) );
  aoim22d1 U5698 ( .A1(n3376), .A2(n3492), .B1(\RegFilePlugin_regFile[12][27] ), .B2(n3377), .Z(n4615) );
  aoim22d1 U5699 ( .A1(n3376), .A2(n3493), .B1(\RegFilePlugin_regFile[12][26] ), .B2(n3375), .Z(n4614) );
  aoim22d1 U5700 ( .A1(n3375), .A2(n3452), .B1(\RegFilePlugin_regFile[12][25] ), .B2(n3377), .Z(n4613) );
  aoim22d1 U5701 ( .A1(n3375), .A2(n3453), .B1(\RegFilePlugin_regFile[12][24] ), .B2(n3376), .Z(n4612) );
  aoim22d1 U5702 ( .A1(n3376), .A2(n3454), .B1(\RegFilePlugin_regFile[12][23] ), .B2(n3377), .Z(n4611) );
  aoim22d1 U5703 ( .A1(n3376), .A2(n3455), .B1(\RegFilePlugin_regFile[12][22] ), .B2(n3376), .Z(n4610) );
  aoim22d1 U5704 ( .A1(n3376), .A2(n3342), .B1(\RegFilePlugin_regFile[12][21] ), .B2(n3376), .Z(n4609) );
  aoim22d1 U5705 ( .A1(n3375), .A2(n3343), .B1(\RegFilePlugin_regFile[12][20] ), .B2(n3377), .Z(n4608) );
  aoim22d1 U5706 ( .A1(n3377), .A2(n3344), .B1(\RegFilePlugin_regFile[12][19] ), .B2(n3376), .Z(n4607) );
  aoim22d1 U5707 ( .A1(n3378), .A2(n3456), .B1(\RegFilePlugin_regFile[12][18] ), .B2(n3376), .Z(n4606) );
  aoim22d1 U5708 ( .A1(n3377), .A2(n3457), .B1(\RegFilePlugin_regFile[12][17] ), .B2(n3377), .Z(n4605) );
  aoim22d1 U5709 ( .A1(n3376), .A2(n3458), .B1(\RegFilePlugin_regFile[12][16] ), .B2(n3377), .Z(n4604) );
  aoim22d1 U5710 ( .A1(n3375), .A2(n3531), .B1(\RegFilePlugin_regFile[12][15] ), .B2(n3377), .Z(n4603) );
  aoim22d1 U5711 ( .A1(n3377), .A2(n3459), .B1(\RegFilePlugin_regFile[12][14] ), .B2(n3377), .Z(n4602) );
  aoim22d1 U5712 ( .A1(n3378), .A2(n3534), .B1(\RegFilePlugin_regFile[12][13] ), .B2(n3377), .Z(n4601) );
  aoim22d1 U5713 ( .A1(n3376), .A2(n3460), .B1(\RegFilePlugin_regFile[12][12] ), .B2(n3377), .Z(n4600) );
  aoim22d1 U5714 ( .A1(n3378), .A2(n3461), .B1(\RegFilePlugin_regFile[12][11] ), .B2(n3376), .Z(n4599) );
  aoim22d1 U5715 ( .A1(n3378), .A2(n3462), .B1(\RegFilePlugin_regFile[12][10] ), .B2(n3375), .Z(n4598) );
  aoim22d1 U5716 ( .A1(n3375), .A2(n3463), .B1(\RegFilePlugin_regFile[12][9] ), 
        .B2(n3378), .Z(n4597) );
  aoim22d1 U5717 ( .A1(n3378), .A2(n3464), .B1(\RegFilePlugin_regFile[12][8] ), 
        .B2(n3375), .Z(n4596) );
  aoim22d1 U5718 ( .A1(n3377), .A2(n3465), .B1(\RegFilePlugin_regFile[12][7] ), 
        .B2(n3375), .Z(n4595) );
  aoim22d1 U5719 ( .A1(n3378), .A2(n3467), .B1(\RegFilePlugin_regFile[12][6] ), 
        .B2(n3375), .Z(n4594) );
  aoim22d1 U5720 ( .A1(n3378), .A2(n3468), .B1(\RegFilePlugin_regFile[12][5] ), 
        .B2(n3378), .Z(n4593) );
  aoim22d1 U5721 ( .A1(n3376), .A2(n3469), .B1(\RegFilePlugin_regFile[12][4] ), 
        .B2(n3378), .Z(n4592) );
  aoim22d1 U5722 ( .A1(n3377), .A2(n3471), .B1(\RegFilePlugin_regFile[12][3] ), 
        .B2(n3378), .Z(n4591) );
  aoim22d1 U5723 ( .A1(n3378), .A2(n3472), .B1(\RegFilePlugin_regFile[12][2] ), 
        .B2(n3378), .Z(n4590) );
  aoim22d1 U5724 ( .A1(n3378), .A2(n3473), .B1(\RegFilePlugin_regFile[12][1] ), 
        .B2(n3378), .Z(n4589) );
  nr02d1 U5725 ( .A1(n3475), .A2(n3392), .ZN(n3379) );
  buffd1 U5726 ( .I(n3379), .Z(n3381) );
  buffd1 U5727 ( .I(n3379), .Z(n3382) );
  aoim22d1 U5728 ( .A1(n3381), .A2(n3482), .B1(\RegFilePlugin_regFile[11][0] ), 
        .B2(n3382), .Z(n4588) );
  buffd1 U5729 ( .I(n3379), .Z(n3380) );
  aoim22d1 U5730 ( .A1(n3380), .A2(n3450), .B1(\RegFilePlugin_regFile[11][31] ), .B2(n3382), .Z(n4587) );
  aoim22d1 U5731 ( .A1(n3381), .A2(n3490), .B1(\RegFilePlugin_regFile[11][30] ), .B2(n3380), .Z(n4586) );
  aoim22d1 U5732 ( .A1(n3381), .A2(n3339), .B1(\RegFilePlugin_regFile[11][29] ), .B2(n3380), .Z(n4585) );
  aoim22d1 U5733 ( .A1(n3379), .A2(n3484), .B1(\RegFilePlugin_regFile[11][28] ), .B2(n3380), .Z(n4584) );
  aoim22d1 U5734 ( .A1(n3381), .A2(n3492), .B1(\RegFilePlugin_regFile[11][27] ), .B2(n3379), .Z(n4583) );
  aoim22d1 U5735 ( .A1(n3381), .A2(n3493), .B1(\RegFilePlugin_regFile[11][26] ), .B2(n3380), .Z(n4582) );
  aoim22d1 U5736 ( .A1(n3380), .A2(n3452), .B1(\RegFilePlugin_regFile[11][25] ), .B2(n3379), .Z(n4581) );
  aoim22d1 U5737 ( .A1(n3380), .A2(n3453), .B1(\RegFilePlugin_regFile[11][24] ), .B2(n3381), .Z(n4580) );
  aoim22d1 U5738 ( .A1(n3381), .A2(n3454), .B1(\RegFilePlugin_regFile[11][23] ), .B2(n3381), .Z(n4579) );
  aoim22d1 U5739 ( .A1(n3381), .A2(n3455), .B1(\RegFilePlugin_regFile[11][22] ), .B2(n3381), .Z(n4578) );
  aoim22d1 U5740 ( .A1(n3381), .A2(n3342), .B1(\RegFilePlugin_regFile[11][21] ), .B2(n3381), .Z(n4577) );
  aoim22d1 U5741 ( .A1(n3380), .A2(n3343), .B1(\RegFilePlugin_regFile[11][20] ), .B2(n3379), .Z(n4576) );
  aoim22d1 U5742 ( .A1(n3379), .A2(n3344), .B1(\RegFilePlugin_regFile[11][19] ), .B2(n3381), .Z(n4575) );
  aoim22d1 U5743 ( .A1(n3382), .A2(n3456), .B1(\RegFilePlugin_regFile[11][18] ), .B2(n3381), .Z(n4574) );
  aoim22d1 U5744 ( .A1(n3379), .A2(n3457), .B1(\RegFilePlugin_regFile[11][17] ), .B2(n3379), .Z(n4573) );
  aoim22d1 U5745 ( .A1(n3381), .A2(n3458), .B1(\RegFilePlugin_regFile[11][16] ), .B2(n3380), .Z(n4572) );
  aoim22d1 U5746 ( .A1(n3380), .A2(n3531), .B1(\RegFilePlugin_regFile[11][15] ), .B2(n3379), .Z(n4571) );
  aoim22d1 U5747 ( .A1(n3379), .A2(n3459), .B1(\RegFilePlugin_regFile[11][14] ), .B2(n3379), .Z(n4570) );
  aoim22d1 U5748 ( .A1(n3382), .A2(n3534), .B1(\RegFilePlugin_regFile[11][13] ), .B2(n3382), .Z(n4569) );
  aoim22d1 U5749 ( .A1(n3381), .A2(n3460), .B1(\RegFilePlugin_regFile[11][12] ), .B2(n3379), .Z(n4568) );
  aoim22d1 U5750 ( .A1(n3382), .A2(n3461), .B1(\RegFilePlugin_regFile[11][11] ), .B2(n3380), .Z(n4567) );
  aoim22d1 U5751 ( .A1(n3382), .A2(n3462), .B1(\RegFilePlugin_regFile[11][10] ), .B2(n3380), .Z(n4566) );
  aoim22d1 U5752 ( .A1(n3380), .A2(n3463), .B1(\RegFilePlugin_regFile[11][9] ), 
        .B2(n3380), .Z(n4565) );
  aoim22d1 U5753 ( .A1(n3382), .A2(n3464), .B1(\RegFilePlugin_regFile[11][8] ), 
        .B2(n3380), .Z(n4564) );
  aoim22d1 U5754 ( .A1(n3379), .A2(n3465), .B1(\RegFilePlugin_regFile[11][7] ), 
        .B2(n3380), .Z(n4563) );
  aoim22d1 U5755 ( .A1(n3382), .A2(n3467), .B1(\RegFilePlugin_regFile[11][6] ), 
        .B2(n3380), .Z(n4562) );
  aoim22d1 U5756 ( .A1(n3382), .A2(n3468), .B1(\RegFilePlugin_regFile[11][5] ), 
        .B2(n3382), .Z(n4561) );
  aoim22d1 U5757 ( .A1(n3381), .A2(n3469), .B1(\RegFilePlugin_regFile[11][4] ), 
        .B2(n3382), .Z(n4560) );
  aoim22d1 U5758 ( .A1(n3379), .A2(n3471), .B1(\RegFilePlugin_regFile[11][3] ), 
        .B2(n3382), .Z(n4559) );
  aoim22d1 U5759 ( .A1(n3382), .A2(n3472), .B1(\RegFilePlugin_regFile[11][2] ), 
        .B2(n3382), .Z(n4558) );
  aoim22d1 U5760 ( .A1(n3382), .A2(n3473), .B1(\RegFilePlugin_regFile[11][1] ), 
        .B2(n3382), .Z(n4557) );
  nr02d1 U5761 ( .A1(n3481), .A2(n3392), .ZN(n3383) );
  buffd1 U5762 ( .I(n3383), .Z(n3384) );
  buffd1 U5763 ( .I(n3383), .Z(n3386) );
  aoim22d1 U5764 ( .A1(n3384), .A2(n3482), .B1(\RegFilePlugin_regFile[10][0] ), 
        .B2(n3386), .Z(n4556) );
  aoim22d1 U5765 ( .A1(n3385), .A2(n3450), .B1(\RegFilePlugin_regFile[10][31] ), .B2(n3386), .Z(n4555) );
  aoim22d1 U5766 ( .A1(n3384), .A2(n3490), .B1(\RegFilePlugin_regFile[10][30] ), .B2(n3383), .Z(n4554) );
  aoim22d1 U5767 ( .A1(n3384), .A2(n3339), .B1(\RegFilePlugin_regFile[10][29] ), .B2(n3383), .Z(n4553) );
  buffd1 U5768 ( .I(n3383), .Z(n3385) );
  aoim22d1 U5769 ( .A1(n3385), .A2(n3476), .B1(\RegFilePlugin_regFile[10][28] ), .B2(n3383), .Z(n4552) );
  aoim22d1 U5770 ( .A1(n3384), .A2(n3492), .B1(\RegFilePlugin_regFile[10][27] ), .B2(n3385), .Z(n4551) );
  aoim22d1 U5771 ( .A1(n3384), .A2(n3493), .B1(\RegFilePlugin_regFile[10][26] ), .B2(n3383), .Z(n4550) );
  aoim22d1 U5772 ( .A1(n3383), .A2(n3452), .B1(\RegFilePlugin_regFile[10][25] ), .B2(n3385), .Z(n4549) );
  aoim22d1 U5773 ( .A1(n3383), .A2(n3453), .B1(\RegFilePlugin_regFile[10][24] ), .B2(n3384), .Z(n4548) );
  aoim22d1 U5774 ( .A1(n3384), .A2(n3454), .B1(\RegFilePlugin_regFile[10][23] ), .B2(n3385), .Z(n4547) );
  aoim22d1 U5775 ( .A1(n3384), .A2(n3455), .B1(\RegFilePlugin_regFile[10][22] ), .B2(n3384), .Z(n4546) );
  aoim22d1 U5776 ( .A1(n3384), .A2(n3342), .B1(\RegFilePlugin_regFile[10][21] ), .B2(n3384), .Z(n4545) );
  aoim22d1 U5777 ( .A1(n3383), .A2(n3343), .B1(\RegFilePlugin_regFile[10][20] ), .B2(n3385), .Z(n4544) );
  aoim22d1 U5778 ( .A1(n3385), .A2(n3344), .B1(\RegFilePlugin_regFile[10][19] ), .B2(n3384), .Z(n4543) );
  aoim22d1 U5779 ( .A1(n3386), .A2(n3456), .B1(\RegFilePlugin_regFile[10][18] ), .B2(n3384), .Z(n4542) );
  aoim22d1 U5780 ( .A1(n3385), .A2(n3457), .B1(\RegFilePlugin_regFile[10][17] ), .B2(n3385), .Z(n4541) );
  aoim22d1 U5781 ( .A1(n3384), .A2(n3458), .B1(\RegFilePlugin_regFile[10][16] ), .B2(n3385), .Z(n4540) );
  aoim22d1 U5782 ( .A1(n3383), .A2(n3531), .B1(\RegFilePlugin_regFile[10][15] ), .B2(n3385), .Z(n4539) );
  aoim22d1 U5783 ( .A1(n3385), .A2(n3459), .B1(\RegFilePlugin_regFile[10][14] ), .B2(n3385), .Z(n4538) );
  aoim22d1 U5784 ( .A1(n3386), .A2(n3534), .B1(\RegFilePlugin_regFile[10][13] ), .B2(n3385), .Z(n4537) );
  aoim22d1 U5785 ( .A1(n3384), .A2(n3460), .B1(\RegFilePlugin_regFile[10][12] ), .B2(n3385), .Z(n4536) );
  aoim22d1 U5786 ( .A1(n3386), .A2(n3461), .B1(\RegFilePlugin_regFile[10][11] ), .B2(n3383), .Z(n4535) );
  aoim22d1 U5787 ( .A1(n3386), .A2(n3462), .B1(\RegFilePlugin_regFile[10][10] ), .B2(n3386), .Z(n4534) );
  aoim22d1 U5788 ( .A1(n3383), .A2(n3463), .B1(\RegFilePlugin_regFile[10][9] ), 
        .B2(n3383), .Z(n4533) );
  aoim22d1 U5789 ( .A1(n3386), .A2(n3464), .B1(\RegFilePlugin_regFile[10][8] ), 
        .B2(n3384), .Z(n4532) );
  aoim22d1 U5790 ( .A1(n3385), .A2(n3465), .B1(\RegFilePlugin_regFile[10][7] ), 
        .B2(n3383), .Z(n4531) );
  aoim22d1 U5791 ( .A1(n3386), .A2(n3467), .B1(\RegFilePlugin_regFile[10][6] ), 
        .B2(n3383), .Z(n4530) );
  aoim22d1 U5792 ( .A1(n3386), .A2(n3468), .B1(\RegFilePlugin_regFile[10][5] ), 
        .B2(n3386), .Z(n4529) );
  aoim22d1 U5793 ( .A1(n3384), .A2(n3469), .B1(\RegFilePlugin_regFile[10][4] ), 
        .B2(n3386), .Z(n4528) );
  aoim22d1 U5794 ( .A1(n3385), .A2(n3471), .B1(\RegFilePlugin_regFile[10][3] ), 
        .B2(n3386), .Z(n4527) );
  aoim22d1 U5795 ( .A1(n3386), .A2(n3472), .B1(\RegFilePlugin_regFile[10][2] ), 
        .B2(n3386), .Z(n4526) );
  aoim22d1 U5796 ( .A1(n3386), .A2(n3473), .B1(\RegFilePlugin_regFile[10][1] ), 
        .B2(n3386), .Z(n4525) );
  nr02d1 U5797 ( .A1(n3489), .A2(n3392), .ZN(n3387) );
  buffd1 U5798 ( .I(n3387), .Z(n3389) );
  buffd1 U5799 ( .I(n3387), .Z(n3390) );
  aoim22d1 U5800 ( .A1(n3389), .A2(n3482), .B1(\RegFilePlugin_regFile[9][0] ), 
        .B2(n3390), .Z(n4524) );
  buffd1 U5801 ( .I(n3387), .Z(n3388) );
  aoim22d1 U5802 ( .A1(n3388), .A2(n3450), .B1(\RegFilePlugin_regFile[9][31] ), 
        .B2(n3390), .Z(n4523) );
  aoim22d1 U5803 ( .A1(n3389), .A2(n3490), .B1(\RegFilePlugin_regFile[9][30] ), 
        .B2(n3388), .Z(n4522) );
  aoim22d1 U5804 ( .A1(n3389), .A2(n3339), .B1(\RegFilePlugin_regFile[9][29] ), 
        .B2(n3388), .Z(n4521) );
  aoim22d1 U5805 ( .A1(n3387), .A2(n3484), .B1(\RegFilePlugin_regFile[9][28] ), 
        .B2(n3388), .Z(n4520) );
  aoim22d1 U5806 ( .A1(n3389), .A2(n3492), .B1(\RegFilePlugin_regFile[9][27] ), 
        .B2(n3390), .Z(n4519) );
  aoim22d1 U5807 ( .A1(n3389), .A2(n3493), .B1(\RegFilePlugin_regFile[9][26] ), 
        .B2(n3388), .Z(n4518) );
  aoim22d1 U5808 ( .A1(n3388), .A2(n3452), .B1(\RegFilePlugin_regFile[9][25] ), 
        .B2(n3389), .Z(n4517) );
  aoim22d1 U5809 ( .A1(n3388), .A2(n3453), .B1(\RegFilePlugin_regFile[9][24] ), 
        .B2(n3389), .Z(n4516) );
  aoim22d1 U5810 ( .A1(n3389), .A2(n3454), .B1(\RegFilePlugin_regFile[9][23] ), 
        .B2(n3387), .Z(n4515) );
  aoim22d1 U5811 ( .A1(n3389), .A2(n3455), .B1(\RegFilePlugin_regFile[9][22] ), 
        .B2(n3389), .Z(n4514) );
  aoim22d1 U5812 ( .A1(n3389), .A2(n3342), .B1(\RegFilePlugin_regFile[9][21] ), 
        .B2(n3389), .Z(n4513) );
  aoim22d1 U5813 ( .A1(n3388), .A2(n3343), .B1(\RegFilePlugin_regFile[9][20] ), 
        .B2(n3387), .Z(n4512) );
  aoim22d1 U5814 ( .A1(n3387), .A2(n3344), .B1(\RegFilePlugin_regFile[9][19] ), 
        .B2(n3389), .Z(n4511) );
  aoim22d1 U5815 ( .A1(n3390), .A2(n3456), .B1(\RegFilePlugin_regFile[9][18] ), 
        .B2(n3389), .Z(n4510) );
  aoim22d1 U5816 ( .A1(n3387), .A2(n3457), .B1(\RegFilePlugin_regFile[9][17] ), 
        .B2(n3387), .Z(n4509) );
  aoim22d1 U5817 ( .A1(n3389), .A2(n3458), .B1(\RegFilePlugin_regFile[9][16] ), 
        .B2(n3387), .Z(n4508) );
  aoim22d1 U5818 ( .A1(n3388), .A2(n3531), .B1(\RegFilePlugin_regFile[9][15] ), 
        .B2(n3387), .Z(n4507) );
  aoim22d1 U5819 ( .A1(n3387), .A2(n3459), .B1(\RegFilePlugin_regFile[9][14] ), 
        .B2(n3387), .Z(n4506) );
  aoim22d1 U5820 ( .A1(n3390), .A2(n3534), .B1(\RegFilePlugin_regFile[9][13] ), 
        .B2(n3388), .Z(n4505) );
  aoim22d1 U5821 ( .A1(n3389), .A2(n3460), .B1(\RegFilePlugin_regFile[9][12] ), 
        .B2(n3387), .Z(n4504) );
  aoim22d1 U5822 ( .A1(n3390), .A2(n3461), .B1(\RegFilePlugin_regFile[9][11] ), 
        .B2(n3388), .Z(n4503) );
  aoim22d1 U5823 ( .A1(n3390), .A2(n3462), .B1(\RegFilePlugin_regFile[9][10] ), 
        .B2(n3388), .Z(n4502) );
  aoim22d1 U5824 ( .A1(n3388), .A2(n3463), .B1(\RegFilePlugin_regFile[9][9] ), 
        .B2(n3388), .Z(n4501) );
  aoim22d1 U5825 ( .A1(n3390), .A2(n3464), .B1(\RegFilePlugin_regFile[9][8] ), 
        .B2(n3388), .Z(n4500) );
  aoim22d1 U5826 ( .A1(n3387), .A2(n3465), .B1(\RegFilePlugin_regFile[9][7] ), 
        .B2(n3388), .Z(n4499) );
  aoim22d1 U5827 ( .A1(n3390), .A2(n3467), .B1(\RegFilePlugin_regFile[9][6] ), 
        .B2(n3388), .Z(n4498) );
  aoim22d1 U5828 ( .A1(n3390), .A2(n3468), .B1(\RegFilePlugin_regFile[9][5] ), 
        .B2(n3390), .Z(n4497) );
  aoim22d1 U5829 ( .A1(n3389), .A2(n3469), .B1(\RegFilePlugin_regFile[9][4] ), 
        .B2(n3390), .Z(n4496) );
  aoim22d1 U5830 ( .A1(n3387), .A2(n3471), .B1(\RegFilePlugin_regFile[9][3] ), 
        .B2(n3390), .Z(n4495) );
  aoim22d1 U5831 ( .A1(n3390), .A2(n3472), .B1(\RegFilePlugin_regFile[9][2] ), 
        .B2(n3390), .Z(n4494) );
  aoim22d1 U5832 ( .A1(n3390), .A2(n3473), .B1(\RegFilePlugin_regFile[9][1] ), 
        .B2(n3390), .Z(n4493) );
  inv0d0 U5833 ( .I(n3391), .ZN(n3393) );
  nr04d0 U5834 ( .A1(_zz_lastStageRegFileWrite_payload_address[9]), .A2(
        _zz_lastStageRegFileWrite_payload_address[8]), .A3(n3393), .A4(n3392), 
        .ZN(n3398) );
  buffd1 U5835 ( .I(n3398), .Z(n3426) );
  buffd1 U5836 ( .I(n3398), .Z(n3425) );
  aoim22d1 U5837 ( .A1(n3426), .A2(n3394), .B1(\RegFilePlugin_regFile[8][0] ), 
        .B2(n3425), .Z(n4492) );
  buffd1 U5838 ( .I(n3398), .Z(n3430) );
  aoim22d1 U5839 ( .A1(n3430), .A2(n3395), .B1(\RegFilePlugin_regFile[8][31] ), 
        .B2(n3426), .Z(n4491) );
  aoim22d1 U5840 ( .A1(n3426), .A2(n3396), .B1(\RegFilePlugin_regFile[8][30] ), 
        .B2(n3425), .Z(n4490) );
  aoim22d1 U5841 ( .A1(n3426), .A2(n3397), .B1(\RegFilePlugin_regFile[8][29] ), 
        .B2(n3425), .Z(n4489) );
  buffd1 U5842 ( .I(n3398), .Z(n3428) );
  aoim22d1 U5843 ( .A1(n3428), .A2(n3399), .B1(\RegFilePlugin_regFile[8][28] ), 
        .B2(n3425), .Z(n4488) );
  aoim22d1 U5844 ( .A1(n3426), .A2(n3400), .B1(\RegFilePlugin_regFile[8][27] ), 
        .B2(n3428), .Z(n4487) );
  aoim22d1 U5845 ( .A1(n3426), .A2(n3401), .B1(\RegFilePlugin_regFile[8][26] ), 
        .B2(n3425), .Z(n4486) );
  aoim22d1 U5846 ( .A1(n3430), .A2(n3402), .B1(\RegFilePlugin_regFile[8][25] ), 
        .B2(n3428), .Z(n4485) );
  aoim22d1 U5847 ( .A1(n3426), .A2(n3403), .B1(\RegFilePlugin_regFile[8][24] ), 
        .B2(n3426), .Z(n4484) );
  aoim22d1 U5848 ( .A1(n3430), .A2(n3404), .B1(\RegFilePlugin_regFile[8][23] ), 
        .B2(n3428), .Z(n4483) );
  aoim22d1 U5849 ( .A1(n3430), .A2(n3405), .B1(\RegFilePlugin_regFile[8][22] ), 
        .B2(n3426), .Z(n4482) );
  aoim22d1 U5850 ( .A1(n3428), .A2(n3406), .B1(\RegFilePlugin_regFile[8][21] ), 
        .B2(n3426), .Z(n4481) );
  aoim22d1 U5851 ( .A1(n3426), .A2(n3407), .B1(\RegFilePlugin_regFile[8][20] ), 
        .B2(n3428), .Z(n4480) );
  aoim22d1 U5852 ( .A1(n3430), .A2(n3408), .B1(\RegFilePlugin_regFile[8][19] ), 
        .B2(n3426), .Z(n4479) );
  aoim22d1 U5853 ( .A1(n3430), .A2(n3409), .B1(\RegFilePlugin_regFile[8][18] ), 
        .B2(n3426), .Z(n4478) );
  aoim22d1 U5854 ( .A1(n3425), .A2(n3410), .B1(\RegFilePlugin_regFile[8][17] ), 
        .B2(n3428), .Z(n4477) );
  aoim22d1 U5855 ( .A1(n3430), .A2(n3411), .B1(\RegFilePlugin_regFile[8][16] ), 
        .B2(n3428), .Z(n4476) );
  aoim22d1 U5856 ( .A1(n3430), .A2(n3412), .B1(\RegFilePlugin_regFile[8][15] ), 
        .B2(n3428), .Z(n4475) );
  aoim22d1 U5857 ( .A1(n3430), .A2(n3413), .B1(\RegFilePlugin_regFile[8][14] ), 
        .B2(n3428), .Z(n4474) );
  aoim22d1 U5858 ( .A1(n3430), .A2(n3414), .B1(\RegFilePlugin_regFile[8][13] ), 
        .B2(n3428), .Z(n4473) );
  aoim22d1 U5859 ( .A1(n3430), .A2(n3415), .B1(\RegFilePlugin_regFile[8][12] ), 
        .B2(n3428), .Z(n4472) );
  aoim22d1 U5860 ( .A1(n3430), .A2(n3416), .B1(\RegFilePlugin_regFile[8][11] ), 
        .B2(n3425), .Z(n4471) );
  aoim22d1 U5861 ( .A1(n3430), .A2(n3417), .B1(\RegFilePlugin_regFile[8][10] ), 
        .B2(n3425), .Z(n4470) );
  aoim22d1 U5862 ( .A1(n3430), .A2(n3418), .B1(\RegFilePlugin_regFile[8][9] ), 
        .B2(n3425), .Z(n4469) );
  aoim22d1 U5863 ( .A1(n3425), .A2(n3419), .B1(\RegFilePlugin_regFile[8][8] ), 
        .B2(n3425), .Z(n4468) );
  aoim22d1 U5864 ( .A1(n3430), .A2(n3420), .B1(\RegFilePlugin_regFile[8][7] ), 
        .B2(n3425), .Z(n4467) );
  aoim22d1 U5865 ( .A1(n3425), .A2(n3421), .B1(\RegFilePlugin_regFile[8][6] ), 
        .B2(n3425), .Z(n4466) );
  aoim22d1 U5866 ( .A1(n3426), .A2(n3422), .B1(\RegFilePlugin_regFile[8][5] ), 
        .B2(n3428), .Z(n4465) );
  aoim22d1 U5867 ( .A1(n3425), .A2(n3423), .B1(\RegFilePlugin_regFile[8][4] ), 
        .B2(n3428), .Z(n4464) );
  aoim22d1 U5868 ( .A1(n3425), .A2(n3424), .B1(\RegFilePlugin_regFile[8][3] ), 
        .B2(n3426), .Z(n4463) );
  aoim22d1 U5869 ( .A1(n3428), .A2(n3427), .B1(\RegFilePlugin_regFile[8][2] ), 
        .B2(n3426), .Z(n4462) );
  aoim22d1 U5870 ( .A1(n3430), .A2(n3429), .B1(\RegFilePlugin_regFile[8][1] ), 
        .B2(n3428), .Z(n4461) );
  nr02d1 U5871 ( .A1(n3434), .A2(n3497), .ZN(n3435) );
  buffd1 U5872 ( .I(n3435), .Z(n3437) );
  buffd1 U5873 ( .I(n3435), .Z(n3438) );
  aoim22d1 U5874 ( .A1(n3437), .A2(n3482), .B1(\RegFilePlugin_regFile[7][0] ), 
        .B2(n3438), .Z(n4460) );
  buffd1 U5875 ( .I(n3435), .Z(n3436) );
  aoim22d1 U5876 ( .A1(n3436), .A2(n3450), .B1(\RegFilePlugin_regFile[7][31] ), 
        .B2(n3438), .Z(n4459) );
  aoim22d1 U5877 ( .A1(n3437), .A2(n3490), .B1(\RegFilePlugin_regFile[7][30] ), 
        .B2(n3436), .Z(n4458) );
  aoim22d1 U5878 ( .A1(n3437), .A2(n3339), .B1(\RegFilePlugin_regFile[7][29] ), 
        .B2(n3436), .Z(n4457) );
  aoim22d1 U5879 ( .A1(n3435), .A2(n3476), .B1(\RegFilePlugin_regFile[7][28] ), 
        .B2(n3436), .Z(n4456) );
  aoim22d1 U5880 ( .A1(n3437), .A2(n3492), .B1(\RegFilePlugin_regFile[7][27] ), 
        .B2(n3435), .Z(n4455) );
  aoim22d1 U5881 ( .A1(n3437), .A2(n3493), .B1(\RegFilePlugin_regFile[7][26] ), 
        .B2(n3436), .Z(n4454) );
  aoim22d1 U5882 ( .A1(n3436), .A2(n3452), .B1(\RegFilePlugin_regFile[7][25] ), 
        .B2(n3438), .Z(n4453) );
  aoim22d1 U5883 ( .A1(n3436), .A2(n3453), .B1(\RegFilePlugin_regFile[7][24] ), 
        .B2(n3437), .Z(n4452) );
  aoim22d1 U5884 ( .A1(n3437), .A2(n3454), .B1(\RegFilePlugin_regFile[7][23] ), 
        .B2(n3437), .Z(n4451) );
  aoim22d1 U5885 ( .A1(n3437), .A2(n3455), .B1(\RegFilePlugin_regFile[7][22] ), 
        .B2(n3437), .Z(n4450) );
  aoim22d1 U5886 ( .A1(n3437), .A2(n3342), .B1(\RegFilePlugin_regFile[7][21] ), 
        .B2(n3437), .Z(n4449) );
  aoim22d1 U5887 ( .A1(n3436), .A2(n3343), .B1(\RegFilePlugin_regFile[7][20] ), 
        .B2(n3435), .Z(n4448) );
  aoim22d1 U5888 ( .A1(n3435), .A2(n3344), .B1(\RegFilePlugin_regFile[7][19] ), 
        .B2(n3437), .Z(n4447) );
  aoim22d1 U5889 ( .A1(n3438), .A2(n3456), .B1(\RegFilePlugin_regFile[7][18] ), 
        .B2(n3437), .Z(n4446) );
  aoim22d1 U5890 ( .A1(n3435), .A2(n3457), .B1(\RegFilePlugin_regFile[7][17] ), 
        .B2(n3435), .Z(n4445) );
  aoim22d1 U5891 ( .A1(n3437), .A2(n3458), .B1(\RegFilePlugin_regFile[7][16] ), 
        .B2(n3435), .Z(n4444) );
  aoim22d1 U5892 ( .A1(n3436), .A2(n3531), .B1(\RegFilePlugin_regFile[7][15] ), 
        .B2(n3435), .Z(n4443) );
  aoim22d1 U5893 ( .A1(n3435), .A2(n3459), .B1(\RegFilePlugin_regFile[7][14] ), 
        .B2(n3435), .Z(n4442) );
  aoim22d1 U5894 ( .A1(n3438), .A2(n3534), .B1(\RegFilePlugin_regFile[7][13] ), 
        .B2(n3435), .Z(n4441) );
  aoim22d1 U5895 ( .A1(n3437), .A2(n3460), .B1(\RegFilePlugin_regFile[7][12] ), 
        .B2(n3435), .Z(n4440) );
  aoim22d1 U5896 ( .A1(n3438), .A2(n3461), .B1(\RegFilePlugin_regFile[7][11] ), 
        .B2(n3436), .Z(n4439) );
  aoim22d1 U5897 ( .A1(n3438), .A2(n3462), .B1(\RegFilePlugin_regFile[7][10] ), 
        .B2(n3436), .Z(n4438) );
  aoim22d1 U5898 ( .A1(n3436), .A2(n3463), .B1(\RegFilePlugin_regFile[7][9] ), 
        .B2(n3436), .Z(n4437) );
  aoim22d1 U5899 ( .A1(n3438), .A2(n3464), .B1(\RegFilePlugin_regFile[7][8] ), 
        .B2(n3436), .Z(n4436) );
  aoim22d1 U5900 ( .A1(n3436), .A2(n3465), .B1(\RegFilePlugin_regFile[7][7] ), 
        .B2(n3436), .Z(n4435) );
  aoim22d1 U5901 ( .A1(n3438), .A2(n3467), .B1(\RegFilePlugin_regFile[7][6] ), 
        .B2(n3436), .Z(n4434) );
  aoim22d1 U5902 ( .A1(n3438), .A2(n3468), .B1(\RegFilePlugin_regFile[7][5] ), 
        .B2(n3438), .Z(n4433) );
  aoim22d1 U5903 ( .A1(n3437), .A2(n3469), .B1(\RegFilePlugin_regFile[7][4] ), 
        .B2(n3438), .Z(n4432) );
  aoim22d1 U5904 ( .A1(n3435), .A2(n3471), .B1(\RegFilePlugin_regFile[7][3] ), 
        .B2(n3438), .Z(n4431) );
  aoim22d1 U5905 ( .A1(n3438), .A2(n3472), .B1(\RegFilePlugin_regFile[7][2] ), 
        .B2(n3438), .Z(n4430) );
  aoim22d1 U5906 ( .A1(n3438), .A2(n3473), .B1(\RegFilePlugin_regFile[7][1] ), 
        .B2(n3438), .Z(n4429) );
  nr02d1 U5907 ( .A1(n3439), .A2(n3497), .ZN(n3440) );
  buffd1 U5908 ( .I(n3440), .Z(n3443) );
  aoim22d1 U5909 ( .A1(n3440), .A2(n3482), .B1(\RegFilePlugin_regFile[6][0] ), 
        .B2(n3443), .Z(n4428) );
  buffd1 U5910 ( .I(n3440), .Z(n3441) );
  aoim22d1 U5911 ( .A1(n3441), .A2(n3450), .B1(\RegFilePlugin_regFile[6][31] ), 
        .B2(n3443), .Z(n4427) );
  aoim22d1 U5912 ( .A1(n3440), .A2(n3490), .B1(\RegFilePlugin_regFile[6][30] ), 
        .B2(n3441), .Z(n4426) );
  aoim22d1 U5913 ( .A1(n3440), .A2(n3339), .B1(\RegFilePlugin_regFile[6][29] ), 
        .B2(n3441), .Z(n4425) );
  buffd1 U5914 ( .I(n3440), .Z(n3442) );
  aoim22d1 U5915 ( .A1(n3442), .A2(n3476), .B1(\RegFilePlugin_regFile[6][28] ), 
        .B2(n3441), .Z(n4424) );
  aoim22d1 U5916 ( .A1(n3440), .A2(n3492), .B1(\RegFilePlugin_regFile[6][27] ), 
        .B2(n3442), .Z(n4423) );
  aoim22d1 U5917 ( .A1(n3440), .A2(n3493), .B1(\RegFilePlugin_regFile[6][26] ), 
        .B2(n3441), .Z(n4422) );
  aoim22d1 U5918 ( .A1(n3441), .A2(n3452), .B1(\RegFilePlugin_regFile[6][25] ), 
        .B2(n3442), .Z(n4421) );
  aoim22d1 U5919 ( .A1(n3441), .A2(n3453), .B1(\RegFilePlugin_regFile[6][24] ), 
        .B2(n3443), .Z(n4420) );
  aoim22d1 U5920 ( .A1(n3440), .A2(n3454), .B1(\RegFilePlugin_regFile[6][23] ), 
        .B2(n3442), .Z(n4419) );
  aoim22d1 U5921 ( .A1(n3440), .A2(n3455), .B1(\RegFilePlugin_regFile[6][22] ), 
        .B2(n3440), .Z(n4418) );
  aoim22d1 U5922 ( .A1(n3441), .A2(n3342), .B1(\RegFilePlugin_regFile[6][21] ), 
        .B2(n3442), .Z(n4417) );
  aoim22d1 U5923 ( .A1(n3441), .A2(n3343), .B1(\RegFilePlugin_regFile[6][20] ), 
        .B2(n3442), .Z(n4416) );
  aoim22d1 U5924 ( .A1(n3442), .A2(n3344), .B1(\RegFilePlugin_regFile[6][19] ), 
        .B2(n3440), .Z(n4415) );
  aoim22d1 U5925 ( .A1(n3443), .A2(n3456), .B1(\RegFilePlugin_regFile[6][18] ), 
        .B2(n3440), .Z(n4414) );
  aoim22d1 U5926 ( .A1(n3442), .A2(n3457), .B1(\RegFilePlugin_regFile[6][17] ), 
        .B2(n3442), .Z(n4413) );
  aoim22d1 U5927 ( .A1(n3440), .A2(n3458), .B1(\RegFilePlugin_regFile[6][16] ), 
        .B2(n3442), .Z(n4412) );
  aoim22d1 U5928 ( .A1(n3441), .A2(n3531), .B1(\RegFilePlugin_regFile[6][15] ), 
        .B2(n3442), .Z(n4411) );
  aoim22d1 U5929 ( .A1(n3442), .A2(n3459), .B1(\RegFilePlugin_regFile[6][14] ), 
        .B2(n3442), .Z(n4410) );
  aoim22d1 U5930 ( .A1(n3443), .A2(n3534), .B1(\RegFilePlugin_regFile[6][13] ), 
        .B2(n3442), .Z(n4409) );
  aoim22d1 U5931 ( .A1(n3440), .A2(n3460), .B1(\RegFilePlugin_regFile[6][12] ), 
        .B2(n3442), .Z(n4408) );
  aoim22d1 U5932 ( .A1(n3443), .A2(n3461), .B1(\RegFilePlugin_regFile[6][11] ), 
        .B2(n3441), .Z(n4407) );
  aoim22d1 U5933 ( .A1(n3443), .A2(n3462), .B1(\RegFilePlugin_regFile[6][10] ), 
        .B2(n3441), .Z(n4406) );
  aoim22d1 U5934 ( .A1(n3441), .A2(n3463), .B1(\RegFilePlugin_regFile[6][9] ), 
        .B2(n3441), .Z(n4405) );
  aoim22d1 U5935 ( .A1(n3443), .A2(n3464), .B1(\RegFilePlugin_regFile[6][8] ), 
        .B2(n3441), .Z(n4404) );
  aoim22d1 U5936 ( .A1(n3442), .A2(n3465), .B1(\RegFilePlugin_regFile[6][7] ), 
        .B2(n3441), .Z(n4403) );
  aoim22d1 U5937 ( .A1(n3443), .A2(n3467), .B1(\RegFilePlugin_regFile[6][6] ), 
        .B2(n3441), .Z(n4402) );
  aoim22d1 U5938 ( .A1(n3443), .A2(n3468), .B1(\RegFilePlugin_regFile[6][5] ), 
        .B2(n3443), .Z(n4401) );
  aoim22d1 U5939 ( .A1(n3440), .A2(n3469), .B1(\RegFilePlugin_regFile[6][4] ), 
        .B2(n3443), .Z(n4400) );
  aoim22d1 U5940 ( .A1(n3442), .A2(n3471), .B1(\RegFilePlugin_regFile[6][3] ), 
        .B2(n3443), .Z(n4399) );
  aoim22d1 U5941 ( .A1(n3443), .A2(n3472), .B1(\RegFilePlugin_regFile[6][2] ), 
        .B2(n3443), .Z(n4398) );
  aoim22d1 U5942 ( .A1(n3443), .A2(n3473), .B1(\RegFilePlugin_regFile[6][1] ), 
        .B2(n3443), .Z(n4397) );
  nr02d1 U5943 ( .A1(n3444), .A2(n3497), .ZN(n3445) );
  buffd1 U5944 ( .I(n3445), .Z(n3447) );
  buffd1 U5945 ( .I(n3445), .Z(n3448) );
  aoim22d1 U5946 ( .A1(n3447), .A2(n3500), .B1(\RegFilePlugin_regFile[5][0] ), 
        .B2(n3448), .Z(n4396) );
  buffd1 U5947 ( .I(n3445), .Z(n3446) );
  aoim22d1 U5948 ( .A1(n3446), .A2(n3450), .B1(\RegFilePlugin_regFile[5][31] ), 
        .B2(n3448), .Z(n4395) );
  aoim22d1 U5949 ( .A1(n3447), .A2(n3490), .B1(\RegFilePlugin_regFile[5][30] ), 
        .B2(n3446), .Z(n4394) );
  aoim22d1 U5950 ( .A1(n3447), .A2(n3339), .B1(\RegFilePlugin_regFile[5][29] ), 
        .B2(n3446), .Z(n4393) );
  aoim22d1 U5951 ( .A1(n3445), .A2(n3476), .B1(\RegFilePlugin_regFile[5][28] ), 
        .B2(n3446), .Z(n4392) );
  aoim22d1 U5952 ( .A1(n3447), .A2(n3492), .B1(\RegFilePlugin_regFile[5][27] ), 
        .B2(n3445), .Z(n4391) );
  aoim22d1 U5953 ( .A1(n3447), .A2(n3493), .B1(\RegFilePlugin_regFile[5][26] ), 
        .B2(n3446), .Z(n4390) );
  aoim22d1 U5954 ( .A1(n3446), .A2(n3452), .B1(\RegFilePlugin_regFile[5][25] ), 
        .B2(n3445), .Z(n4389) );
  aoim22d1 U5955 ( .A1(n3446), .A2(n3453), .B1(\RegFilePlugin_regFile[5][24] ), 
        .B2(n3447), .Z(n4388) );
  aoim22d1 U5956 ( .A1(n3447), .A2(n3454), .B1(\RegFilePlugin_regFile[5][23] ), 
        .B2(n3447), .Z(n4387) );
  aoim22d1 U5957 ( .A1(n3447), .A2(n3455), .B1(\RegFilePlugin_regFile[5][22] ), 
        .B2(n3447), .Z(n4386) );
  aoim22d1 U5958 ( .A1(n3447), .A2(n3342), .B1(\RegFilePlugin_regFile[5][21] ), 
        .B2(n3447), .Z(n4385) );
  aoim22d1 U5959 ( .A1(n3446), .A2(n3521), .B1(\RegFilePlugin_regFile[5][20] ), 
        .B2(n3445), .Z(n4384) );
  aoim22d1 U5960 ( .A1(n3445), .A2(n3344), .B1(\RegFilePlugin_regFile[5][19] ), 
        .B2(n3447), .Z(n4383) );
  aoim22d1 U5961 ( .A1(n3448), .A2(n3456), .B1(\RegFilePlugin_regFile[5][18] ), 
        .B2(n3447), .Z(n4382) );
  aoim22d1 U5962 ( .A1(n3445), .A2(n3457), .B1(\RegFilePlugin_regFile[5][17] ), 
        .B2(n3445), .Z(n4381) );
  aoim22d1 U5963 ( .A1(n3447), .A2(n3458), .B1(\RegFilePlugin_regFile[5][16] ), 
        .B2(n3445), .Z(n4380) );
  aoim22d1 U5964 ( .A1(n3446), .A2(n3531), .B1(\RegFilePlugin_regFile[5][15] ), 
        .B2(n3446), .Z(n4379) );
  aoim22d1 U5965 ( .A1(n3445), .A2(n3459), .B1(\RegFilePlugin_regFile[5][14] ), 
        .B2(n3445), .Z(n4378) );
  aoim22d1 U5966 ( .A1(n3448), .A2(n3534), .B1(\RegFilePlugin_regFile[5][13] ), 
        .B2(n3445), .Z(n4377) );
  aoim22d1 U5967 ( .A1(n3447), .A2(n3460), .B1(\RegFilePlugin_regFile[5][12] ), 
        .B2(n3445), .Z(n4376) );
  aoim22d1 U5968 ( .A1(n3448), .A2(n3461), .B1(\RegFilePlugin_regFile[5][11] ), 
        .B2(n3446), .Z(n4375) );
  aoim22d1 U5969 ( .A1(n3448), .A2(n3462), .B1(\RegFilePlugin_regFile[5][10] ), 
        .B2(n3446), .Z(n4374) );
  aoim22d1 U5970 ( .A1(n3446), .A2(n3463), .B1(\RegFilePlugin_regFile[5][9] ), 
        .B2(n3446), .Z(n4373) );
  aoim22d1 U5971 ( .A1(n3448), .A2(n3464), .B1(\RegFilePlugin_regFile[5][8] ), 
        .B2(n3446), .Z(n4372) );
  aoim22d1 U5972 ( .A1(n3448), .A2(n3465), .B1(\RegFilePlugin_regFile[5][7] ), 
        .B2(n3446), .Z(n4371) );
  aoim22d1 U5973 ( .A1(n3448), .A2(n3467), .B1(\RegFilePlugin_regFile[5][6] ), 
        .B2(n3446), .Z(n4370) );
  aoim22d1 U5974 ( .A1(n3448), .A2(n3468), .B1(\RegFilePlugin_regFile[5][5] ), 
        .B2(n3448), .Z(n4369) );
  aoim22d1 U5975 ( .A1(n3447), .A2(n3469), .B1(\RegFilePlugin_regFile[5][4] ), 
        .B2(n3448), .Z(n4368) );
  aoim22d1 U5976 ( .A1(n3445), .A2(n3471), .B1(\RegFilePlugin_regFile[5][3] ), 
        .B2(n3448), .Z(n4367) );
  aoim22d1 U5977 ( .A1(n3448), .A2(n3472), .B1(\RegFilePlugin_regFile[5][2] ), 
        .B2(n3448), .Z(n4366) );
  aoim22d1 U5978 ( .A1(n3448), .A2(n3473), .B1(\RegFilePlugin_regFile[5][1] ), 
        .B2(n3448), .Z(n4365) );
  nr02d1 U5979 ( .A1(n3449), .A2(n3497), .ZN(n3451) );
  buffd1 U5980 ( .I(n3451), .Z(n3470) );
  buffd1 U5981 ( .I(n3451), .Z(n3474) );
  aoim22d1 U5982 ( .A1(n3470), .A2(n3500), .B1(\RegFilePlugin_regFile[4][0] ), 
        .B2(n3474), .Z(n4364) );
  buffd1 U5983 ( .I(n3451), .Z(n3466) );
  aoim22d1 U5984 ( .A1(n3466), .A2(n3450), .B1(\RegFilePlugin_regFile[4][31] ), 
        .B2(n3474), .Z(n4363) );
  aoim22d1 U5985 ( .A1(n3470), .A2(n3490), .B1(\RegFilePlugin_regFile[4][30] ), 
        .B2(n3466), .Z(n4362) );
  aoim22d1 U5986 ( .A1(n3470), .A2(n3339), .B1(\RegFilePlugin_regFile[4][29] ), 
        .B2(n3466), .Z(n4361) );
  aoim22d1 U5987 ( .A1(n3451), .A2(n3476), .B1(\RegFilePlugin_regFile[4][28] ), 
        .B2(n3466), .Z(n4360) );
  aoim22d1 U5988 ( .A1(n3470), .A2(n3492), .B1(\RegFilePlugin_regFile[4][27] ), 
        .B2(n3466), .Z(n4359) );
  aoim22d1 U5989 ( .A1(n3470), .A2(n3493), .B1(\RegFilePlugin_regFile[4][26] ), 
        .B2(n3466), .Z(n4358) );
  aoim22d1 U5990 ( .A1(n3466), .A2(n3452), .B1(\RegFilePlugin_regFile[4][25] ), 
        .B2(n3451), .Z(n4357) );
  aoim22d1 U5991 ( .A1(n3466), .A2(n3453), .B1(\RegFilePlugin_regFile[4][24] ), 
        .B2(n3470), .Z(n4356) );
  aoim22d1 U5992 ( .A1(n3470), .A2(n3454), .B1(\RegFilePlugin_regFile[4][23] ), 
        .B2(n3451), .Z(n4355) );
  aoim22d1 U5993 ( .A1(n3470), .A2(n3455), .B1(\RegFilePlugin_regFile[4][22] ), 
        .B2(n3470), .Z(n4354) );
  aoim22d1 U5994 ( .A1(n3470), .A2(n3342), .B1(\RegFilePlugin_regFile[4][21] ), 
        .B2(n3470), .Z(n4353) );
  aoim22d1 U5995 ( .A1(n3466), .A2(n3343), .B1(\RegFilePlugin_regFile[4][20] ), 
        .B2(n3451), .Z(n4352) );
  aoim22d1 U5996 ( .A1(n3474), .A2(n3344), .B1(\RegFilePlugin_regFile[4][19] ), 
        .B2(n3470), .Z(n4351) );
  aoim22d1 U5997 ( .A1(n3474), .A2(n3456), .B1(\RegFilePlugin_regFile[4][18] ), 
        .B2(n3470), .Z(n4350) );
  aoim22d1 U5998 ( .A1(n3451), .A2(n3457), .B1(\RegFilePlugin_regFile[4][17] ), 
        .B2(n3451), .Z(n4349) );
  aoim22d1 U5999 ( .A1(n3470), .A2(n3458), .B1(\RegFilePlugin_regFile[4][16] ), 
        .B2(n3470), .Z(n4348) );
  aoim22d1 U6000 ( .A1(n3466), .A2(n3531), .B1(\RegFilePlugin_regFile[4][15] ), 
        .B2(n3451), .Z(n4347) );
  aoim22d1 U6001 ( .A1(n3451), .A2(n3459), .B1(\RegFilePlugin_regFile[4][14] ), 
        .B2(n3451), .Z(n4346) );
  aoim22d1 U6002 ( .A1(n3474), .A2(n3534), .B1(\RegFilePlugin_regFile[4][13] ), 
        .B2(n3451), .Z(n4345) );
  aoim22d1 U6003 ( .A1(n3470), .A2(n3460), .B1(\RegFilePlugin_regFile[4][12] ), 
        .B2(n3451), .Z(n4344) );
  aoim22d1 U6004 ( .A1(n3474), .A2(n3461), .B1(\RegFilePlugin_regFile[4][11] ), 
        .B2(n3466), .Z(n4343) );
  aoim22d1 U6005 ( .A1(n3474), .A2(n3462), .B1(\RegFilePlugin_regFile[4][10] ), 
        .B2(n3466), .Z(n4342) );
  aoim22d1 U6006 ( .A1(n3466), .A2(n3463), .B1(\RegFilePlugin_regFile[4][9] ), 
        .B2(n3466), .Z(n4341) );
  aoim22d1 U6007 ( .A1(n3474), .A2(n3464), .B1(\RegFilePlugin_regFile[4][8] ), 
        .B2(n3466), .Z(n4340) );
  aoim22d1 U6008 ( .A1(n3451), .A2(n3465), .B1(\RegFilePlugin_regFile[4][7] ), 
        .B2(n3466), .Z(n4339) );
  aoim22d1 U6009 ( .A1(n3474), .A2(n3467), .B1(\RegFilePlugin_regFile[4][6] ), 
        .B2(n3466), .Z(n4338) );
  aoim22d1 U6010 ( .A1(n3474), .A2(n3468), .B1(\RegFilePlugin_regFile[4][5] ), 
        .B2(n3474), .Z(n4337) );
  aoim22d1 U6011 ( .A1(n3470), .A2(n3469), .B1(\RegFilePlugin_regFile[4][4] ), 
        .B2(n3474), .Z(n4336) );
  aoim22d1 U6012 ( .A1(n3451), .A2(n3471), .B1(\RegFilePlugin_regFile[4][3] ), 
        .B2(n3474), .Z(n4335) );
  aoim22d1 U6013 ( .A1(n3474), .A2(n3472), .B1(\RegFilePlugin_regFile[4][2] ), 
        .B2(n3474), .Z(n4334) );
  aoim22d1 U6014 ( .A1(n3474), .A2(n3473), .B1(\RegFilePlugin_regFile[4][1] ), 
        .B2(n3474), .Z(n4333) );
  nr02d1 U6015 ( .A1(n3475), .A2(n3497), .ZN(n3477) );
  buffd1 U6016 ( .I(n3477), .Z(n3478) );
  buffd1 U6017 ( .I(n3477), .Z(n3480) );
  aoim22d1 U6018 ( .A1(n3478), .A2(n3482), .B1(\RegFilePlugin_regFile[3][0] ), 
        .B2(n3480), .Z(n4332) );
  buffd1 U6019 ( .I(n3477), .Z(n3479) );
  aoim22d1 U6020 ( .A1(n3479), .A2(n3338), .B1(\RegFilePlugin_regFile[3][31] ), 
        .B2(n3480), .Z(n4331) );
  aoim22d1 U6021 ( .A1(n3478), .A2(n3490), .B1(\RegFilePlugin_regFile[3][30] ), 
        .B2(n3479), .Z(n4330) );
  aoim22d1 U6022 ( .A1(n3478), .A2(n3505), .B1(\RegFilePlugin_regFile[3][29] ), 
        .B2(n3479), .Z(n4329) );
  aoim22d1 U6023 ( .A1(n3480), .A2(n3476), .B1(\RegFilePlugin_regFile[3][28] ), 
        .B2(n3479), .Z(n4328) );
  aoim22d1 U6024 ( .A1(n3478), .A2(n3492), .B1(\RegFilePlugin_regFile[3][27] ), 
        .B2(n3477), .Z(n4327) );
  aoim22d1 U6025 ( .A1(n3478), .A2(n3493), .B1(\RegFilePlugin_regFile[3][26] ), 
        .B2(n3479), .Z(n4326) );
  aoim22d1 U6026 ( .A1(n3478), .A2(n3512), .B1(\RegFilePlugin_regFile[3][25] ), 
        .B2(n3477), .Z(n4325) );
  aoim22d1 U6027 ( .A1(n3479), .A2(n3341), .B1(\RegFilePlugin_regFile[3][24] ), 
        .B2(n3478), .Z(n4324) );
  aoim22d1 U6028 ( .A1(n3478), .A2(n3454), .B1(\RegFilePlugin_regFile[3][23] ), 
        .B2(n3478), .Z(n4323) );
  aoim22d1 U6029 ( .A1(n3480), .A2(n3517), .B1(\RegFilePlugin_regFile[3][22] ), 
        .B2(n3478), .Z(n4322) );
  aoim22d1 U6030 ( .A1(n3479), .A2(n3519), .B1(\RegFilePlugin_regFile[3][21] ), 
        .B2(n3478), .Z(n4321) );
  aoim22d1 U6031 ( .A1(n3479), .A2(n3521), .B1(\RegFilePlugin_regFile[3][20] ), 
        .B2(n3477), .Z(n4320) );
  aoim22d1 U6032 ( .A1(n3478), .A2(n3523), .B1(\RegFilePlugin_regFile[3][19] ), 
        .B2(n3478), .Z(n4319) );
  aoim22d1 U6033 ( .A1(n3480), .A2(n3456), .B1(\RegFilePlugin_regFile[3][18] ), 
        .B2(n3478), .Z(n4318) );
  aoim22d1 U6034 ( .A1(n3477), .A2(n3527), .B1(\RegFilePlugin_regFile[3][17] ), 
        .B2(n3477), .Z(n4317) );
  aoim22d1 U6035 ( .A1(n3480), .A2(n3529), .B1(\RegFilePlugin_regFile[3][16] ), 
        .B2(n3477), .Z(n4316) );
  aoim22d1 U6036 ( .A1(n3480), .A2(n3531), .B1(\RegFilePlugin_regFile[3][15] ), 
        .B2(n3477), .Z(n4315) );
  aoim22d1 U6037 ( .A1(n3480), .A2(n3459), .B1(\RegFilePlugin_regFile[3][14] ), 
        .B2(n3477), .Z(n4314) );
  aoim22d1 U6038 ( .A1(n3480), .A2(n3534), .B1(\RegFilePlugin_regFile[3][13] ), 
        .B2(n3477), .Z(n4313) );
  aoim22d1 U6039 ( .A1(n3480), .A2(n3460), .B1(\RegFilePlugin_regFile[3][12] ), 
        .B2(n3477), .Z(n4312) );
  aoim22d1 U6040 ( .A1(n3479), .A2(n3461), .B1(\RegFilePlugin_regFile[3][11] ), 
        .B2(n3479), .Z(n4311) );
  aoim22d1 U6041 ( .A1(n3479), .A2(n3462), .B1(\RegFilePlugin_regFile[3][10] ), 
        .B2(n3479), .Z(n4310) );
  aoim22d1 U6042 ( .A1(n3478), .A2(n3463), .B1(\RegFilePlugin_regFile[3][9] ), 
        .B2(n3479), .Z(n4309) );
  aoim22d1 U6043 ( .A1(n3477), .A2(n3541), .B1(\RegFilePlugin_regFile[3][8] ), 
        .B2(n3479), .Z(n4308) );
  aoim22d1 U6044 ( .A1(n3480), .A2(n3543), .B1(\RegFilePlugin_regFile[3][7] ), 
        .B2(n3479), .Z(n4307) );
  aoim22d1 U6045 ( .A1(n3478), .A2(n3467), .B1(\RegFilePlugin_regFile[3][6] ), 
        .B2(n3479), .Z(n4306) );
  aoim22d1 U6046 ( .A1(n3478), .A2(n3468), .B1(\RegFilePlugin_regFile[3][5] ), 
        .B2(n3480), .Z(n4305) );
  aoim22d1 U6047 ( .A1(n3477), .A2(n3469), .B1(\RegFilePlugin_regFile[3][4] ), 
        .B2(n3480), .Z(n4304) );
  aoim22d1 U6048 ( .A1(n3479), .A2(n3551), .B1(\RegFilePlugin_regFile[3][3] ), 
        .B2(n3480), .Z(n4303) );
  aoim22d1 U6049 ( .A1(n3477), .A2(n3472), .B1(\RegFilePlugin_regFile[3][2] ), 
        .B2(n3480), .Z(n4302) );
  aoim22d1 U6050 ( .A1(n3480), .A2(n3554), .B1(\RegFilePlugin_regFile[3][1] ), 
        .B2(n3480), .Z(n4301) );
  nr02d1 U6051 ( .A1(n3481), .A2(n3497), .ZN(n3483) );
  buffd1 U6052 ( .I(n3483), .Z(n3486) );
  buffd1 U6053 ( .I(n3483), .Z(n3488) );
  aoim22d1 U6054 ( .A1(n3486), .A2(n3482), .B1(\RegFilePlugin_regFile[2][0] ), 
        .B2(n3488), .Z(n4300) );
  buffd1 U6055 ( .I(n3483), .Z(n3487) );
  aoim22d1 U6056 ( .A1(n3487), .A2(n3338), .B1(\RegFilePlugin_regFile[2][31] ), 
        .B2(n3488), .Z(n4299) );
  aoim22d1 U6057 ( .A1(n3486), .A2(n3490), .B1(\RegFilePlugin_regFile[2][30] ), 
        .B2(n3483), .Z(n4298) );
  aoim22d1 U6058 ( .A1(n3486), .A2(n3505), .B1(\RegFilePlugin_regFile[2][29] ), 
        .B2(n3483), .Z(n4297) );
  aoim22d1 U6059 ( .A1(n3486), .A2(n3484), .B1(\RegFilePlugin_regFile[2][28] ), 
        .B2(n3483), .Z(n4296) );
  aoim22d1 U6060 ( .A1(n3486), .A2(n3492), .B1(\RegFilePlugin_regFile[2][27] ), 
        .B2(n3487), .Z(n4295) );
  aoim22d1 U6061 ( .A1(n3486), .A2(n3493), .B1(\RegFilePlugin_regFile[2][26] ), 
        .B2(n3483), .Z(n4294) );
  aoim22d1 U6062 ( .A1(n3483), .A2(n3512), .B1(\RegFilePlugin_regFile[2][25] ), 
        .B2(n3487), .Z(n4293) );
  aoim22d1 U6063 ( .A1(n3487), .A2(n3453), .B1(\RegFilePlugin_regFile[2][24] ), 
        .B2(n3486), .Z(n4292) );
  aoim22d1 U6064 ( .A1(n3486), .A2(n3454), .B1(\RegFilePlugin_regFile[2][23] ), 
        .B2(n3487), .Z(n4291) );
  aoim22d1 U6065 ( .A1(n3487), .A2(n3517), .B1(\RegFilePlugin_regFile[2][22] ), 
        .B2(n3486), .Z(n4290) );
  aoim22d1 U6066 ( .A1(n3487), .A2(n3519), .B1(\RegFilePlugin_regFile[2][21] ), 
        .B2(n3486), .Z(n4289) );
  aoim22d1 U6067 ( .A1(n3486), .A2(n3521), .B1(\RegFilePlugin_regFile[2][20] ), 
        .B2(n3487), .Z(n4288) );
  aoim22d1 U6068 ( .A1(n3483), .A2(n3523), .B1(\RegFilePlugin_regFile[2][19] ), 
        .B2(n3486), .Z(n4287) );
  aoim22d1 U6069 ( .A1(n3488), .A2(n3456), .B1(\RegFilePlugin_regFile[2][18] ), 
        .B2(n3486), .Z(n4286) );
  aoim22d1 U6070 ( .A1(n3488), .A2(n3527), .B1(\RegFilePlugin_regFile[2][17] ), 
        .B2(n3487), .Z(n4285) );
  aoim22d1 U6071 ( .A1(n3488), .A2(n3529), .B1(\RegFilePlugin_regFile[2][16] ), 
        .B2(n3487), .Z(n4284) );
  aoim22d1 U6072 ( .A1(n3488), .A2(n3531), .B1(\RegFilePlugin_regFile[2][15] ), 
        .B2(n3487), .Z(n4283) );
  aoim22d1 U6073 ( .A1(n3488), .A2(n3459), .B1(\RegFilePlugin_regFile[2][14] ), 
        .B2(n3487), .Z(n4282) );
  aoim22d1 U6074 ( .A1(n3488), .A2(n3485), .B1(\RegFilePlugin_regFile[2][13] ), 
        .B2(n3487), .Z(n4281) );
  aoim22d1 U6075 ( .A1(n3488), .A2(n3460), .B1(\RegFilePlugin_regFile[2][12] ), 
        .B2(n3487), .Z(n4280) );
  aoim22d1 U6076 ( .A1(n3488), .A2(n3461), .B1(\RegFilePlugin_regFile[2][11] ), 
        .B2(n3483), .Z(n4279) );
  aoim22d1 U6077 ( .A1(n3487), .A2(n3462), .B1(\RegFilePlugin_regFile[2][10] ), 
        .B2(n3483), .Z(n4278) );
  aoim22d1 U6078 ( .A1(n3486), .A2(n3463), .B1(\RegFilePlugin_regFile[2][9] ), 
        .B2(n3486), .Z(n4277) );
  aoim22d1 U6079 ( .A1(n3483), .A2(n3541), .B1(\RegFilePlugin_regFile[2][8] ), 
        .B2(n3483), .Z(n4276) );
  aoim22d1 U6080 ( .A1(n3488), .A2(n3543), .B1(\RegFilePlugin_regFile[2][7] ), 
        .B2(n3487), .Z(n4275) );
  aoim22d1 U6081 ( .A1(n3486), .A2(n3467), .B1(\RegFilePlugin_regFile[2][6] ), 
        .B2(n3483), .Z(n4274) );
  aoim22d1 U6082 ( .A1(n3486), .A2(n3468), .B1(\RegFilePlugin_regFile[2][5] ), 
        .B2(n3488), .Z(n4273) );
  aoim22d1 U6083 ( .A1(n3483), .A2(n3469), .B1(\RegFilePlugin_regFile[2][4] ), 
        .B2(n3488), .Z(n4272) );
  aoim22d1 U6084 ( .A1(n3487), .A2(n3551), .B1(\RegFilePlugin_regFile[2][3] ), 
        .B2(n3488), .Z(n4271) );
  aoim22d1 U6085 ( .A1(n3483), .A2(n3472), .B1(\RegFilePlugin_regFile[2][2] ), 
        .B2(n3488), .Z(n4270) );
  aoim22d1 U6086 ( .A1(n3488), .A2(n3554), .B1(\RegFilePlugin_regFile[2][1] ), 
        .B2(n3488), .Z(n4269) );
  nr02d1 U6087 ( .A1(n3489), .A2(n3497), .ZN(n3491) );
  buffd1 U6088 ( .I(n3491), .Z(n3494) );
  aoim22d1 U6089 ( .A1(n3494), .A2(n3500), .B1(\RegFilePlugin_regFile[1][0] ), 
        .B2(n3494), .Z(n4268) );
  aoim22d1 U6090 ( .A1(n3491), .A2(n3338), .B1(\RegFilePlugin_regFile[1][31] ), 
        .B2(n3491), .Z(n4267) );
  buffd1 U6091 ( .I(n3491), .Z(n3496) );
  aoim22d1 U6092 ( .A1(n3494), .A2(n3490), .B1(\RegFilePlugin_regFile[1][30] ), 
        .B2(n3496), .Z(n4266) );
  aoim22d1 U6093 ( .A1(n3494), .A2(n3505), .B1(\RegFilePlugin_regFile[1][29] ), 
        .B2(n3496), .Z(n4265) );
  aoim22d1 U6094 ( .A1(n3496), .A2(n3476), .B1(\RegFilePlugin_regFile[1][28] ), 
        .B2(n3496), .Z(n4264) );
  buffd1 U6095 ( .I(n3491), .Z(n3495) );
  aoim22d1 U6096 ( .A1(n3494), .A2(n3492), .B1(\RegFilePlugin_regFile[1][27] ), 
        .B2(n3495), .Z(n4263) );
  aoim22d1 U6097 ( .A1(n3494), .A2(n3493), .B1(\RegFilePlugin_regFile[1][26] ), 
        .B2(n3496), .Z(n4262) );
  aoim22d1 U6098 ( .A1(n3494), .A2(n3512), .B1(\RegFilePlugin_regFile[1][25] ), 
        .B2(n3495), .Z(n4261) );
  aoim22d1 U6099 ( .A1(n3496), .A2(n3341), .B1(\RegFilePlugin_regFile[1][24] ), 
        .B2(n3494), .Z(n4260) );
  aoim22d1 U6100 ( .A1(n3494), .A2(n3454), .B1(\RegFilePlugin_regFile[1][23] ), 
        .B2(n3495), .Z(n4259) );
  aoim22d1 U6101 ( .A1(n3491), .A2(n3517), .B1(\RegFilePlugin_regFile[1][22] ), 
        .B2(n3494), .Z(n4258) );
  aoim22d1 U6102 ( .A1(n3495), .A2(n3519), .B1(\RegFilePlugin_regFile[1][21] ), 
        .B2(n3494), .Z(n4257) );
  aoim22d1 U6103 ( .A1(n3495), .A2(n3521), .B1(\RegFilePlugin_regFile[1][20] ), 
        .B2(n3495), .Z(n4256) );
  aoim22d1 U6104 ( .A1(n3494), .A2(n3523), .B1(\RegFilePlugin_regFile[1][19] ), 
        .B2(n3494), .Z(n4255) );
  aoim22d1 U6105 ( .A1(n3495), .A2(n3456), .B1(\RegFilePlugin_regFile[1][18] ), 
        .B2(n3494), .Z(n4254) );
  aoim22d1 U6106 ( .A1(n3496), .A2(n3527), .B1(\RegFilePlugin_regFile[1][17] ), 
        .B2(n3495), .Z(n4253) );
  aoim22d1 U6107 ( .A1(n3491), .A2(n3529), .B1(\RegFilePlugin_regFile[1][16] ), 
        .B2(n3495), .Z(n4252) );
  aoim22d1 U6108 ( .A1(n3491), .A2(n3531), .B1(\RegFilePlugin_regFile[1][15] ), 
        .B2(n3495), .Z(n4251) );
  aoim22d1 U6109 ( .A1(n3491), .A2(n3459), .B1(\RegFilePlugin_regFile[1][14] ), 
        .B2(n3495), .Z(n4250) );
  aoim22d1 U6110 ( .A1(n3496), .A2(n3534), .B1(\RegFilePlugin_regFile[1][13] ), 
        .B2(n3495), .Z(n4249) );
  aoim22d1 U6111 ( .A1(n3491), .A2(n3460), .B1(\RegFilePlugin_regFile[1][12] ), 
        .B2(n3495), .Z(n4248) );
  aoim22d1 U6112 ( .A1(n3495), .A2(n3461), .B1(\RegFilePlugin_regFile[1][11] ), 
        .B2(n3496), .Z(n4247) );
  aoim22d1 U6113 ( .A1(n3495), .A2(n3462), .B1(\RegFilePlugin_regFile[1][10] ), 
        .B2(n3496), .Z(n4246) );
  aoim22d1 U6114 ( .A1(n3494), .A2(n3463), .B1(\RegFilePlugin_regFile[1][9] ), 
        .B2(n3496), .Z(n4245) );
  aoim22d1 U6115 ( .A1(n3494), .A2(n3541), .B1(\RegFilePlugin_regFile[1][8] ), 
        .B2(n3496), .Z(n4244) );
  aoim22d1 U6116 ( .A1(n3495), .A2(n3543), .B1(\RegFilePlugin_regFile[1][7] ), 
        .B2(n3496), .Z(n4243) );
  aoim22d1 U6117 ( .A1(n3496), .A2(n3467), .B1(\RegFilePlugin_regFile[1][6] ), 
        .B2(n3496), .Z(n4242) );
  aoim22d1 U6118 ( .A1(n3494), .A2(n3468), .B1(\RegFilePlugin_regFile[1][5] ), 
        .B2(n3491), .Z(n4241) );
  aoim22d1 U6119 ( .A1(n3496), .A2(n3469), .B1(\RegFilePlugin_regFile[1][4] ), 
        .B2(n3491), .Z(n4240) );
  aoim22d1 U6120 ( .A1(n3495), .A2(n3551), .B1(\RegFilePlugin_regFile[1][3] ), 
        .B2(n3491), .Z(n4239) );
  aoim22d1 U6121 ( .A1(n3496), .A2(n3472), .B1(\RegFilePlugin_regFile[1][2] ), 
        .B2(n3491), .Z(n4238) );
  aoim22d1 U6122 ( .A1(n3491), .A2(n3554), .B1(\RegFilePlugin_regFile[1][1] ), 
        .B2(n3491), .Z(n4237) );
  inv0d0 U6123 ( .I(\RegFilePlugin_regFile[0][0] ), .ZN(n3501) );
  or02d1 U6124 ( .A1(n3498), .A2(n3497), .Z(n3555) );
  buffd1 U6125 ( .I(n3555), .Z(n3549) );
  nd02d1 U6126 ( .A1(n3499), .A2(n3549), .ZN(n3545) );
  buffd1 U6127 ( .I(n3545), .Z(n3556) );
  aoi22d1 U6128 ( .A1(n3501), .A2(n3555), .B1(n3556), .B2(n3500), .ZN(n4236)
         );
  mx02d1 U6129 ( .I0(execute_RS1[0]), .I1(_zz_RegFilePlugin_regFile_port0[0]), 
        .S(n3516), .Z(n4235) );
  inv0d0 U6130 ( .I(\RegFilePlugin_regFile[0][31] ), .ZN(n3502) );
  oai22d1 U6131 ( .A1(n3502), .A2(n3545), .B1(n3338), .B2(n3549), .ZN(n4234)
         );
  mx02d1 U6132 ( .I0(execute_RS1[31]), .I1(_zz_RegFilePlugin_regFile_port0[31]), .S(n3526), .Z(n4233) );
  mx02d1 U6133 ( .I0(execute_RS2[31]), .I1(_zz_RegFilePlugin_regFile_port1[31]), .S(n3516), .Z(n4232) );
  inv0d0 U6134 ( .I(\RegFilePlugin_regFile[0][30] ), .ZN(n3504) );
  aoi22d1 U6135 ( .A1(n3504), .A2(n3549), .B1(n3503), .B2(n3545), .ZN(n4231)
         );
  mx02d1 U6136 ( .I0(execute_RS1[30]), .I1(_zz_RegFilePlugin_regFile_port0[30]), .S(n3516), .Z(n4230) );
  mx02d1 U6137 ( .I0(execute_RS2[30]), .I1(_zz_RegFilePlugin_regFile_port1[30]), .S(n3516), .Z(n4229) );
  inv0d0 U6138 ( .I(\RegFilePlugin_regFile[0][29] ), .ZN(n3506) );
  oai22d1 U6139 ( .A1(n3506), .A2(n3556), .B1(n3505), .B2(n3549), .ZN(n4228)
         );
  mx02d1 U6140 ( .I0(execute_RS1[29]), .I1(_zz_RegFilePlugin_regFile_port0[29]), .S(n3516), .Z(n4227) );
  mx02d1 U6141 ( .I0(execute_RS2[29]), .I1(_zz_RegFilePlugin_regFile_port1[29]), .S(n3516), .Z(n4226) );
  inv0d0 U6142 ( .I(\RegFilePlugin_regFile[0][28] ), .ZN(n3507) );
  aoi22d1 U6143 ( .A1(n3507), .A2(n3555), .B1(n3484), .B2(n3545), .ZN(n4225)
         );
  mx02d1 U6144 ( .I0(execute_RS1[28]), .I1(_zz_RegFilePlugin_regFile_port0[28]), .S(n3516), .Z(n4224) );
  mx02d1 U6145 ( .I0(execute_RS2[28]), .I1(_zz_RegFilePlugin_regFile_port1[28]), .S(n3516), .Z(n4223) );
  inv0d0 U6146 ( .I(\RegFilePlugin_regFile[0][27] ), .ZN(n3509) );
  aoi22d1 U6147 ( .A1(n3509), .A2(n3555), .B1(n3508), .B2(n3545), .ZN(n4222)
         );
  mx02d1 U6148 ( .I0(execute_RS1[27]), .I1(_zz_RegFilePlugin_regFile_port0[27]), .S(n3516), .Z(n4221) );
  mx02d1 U6149 ( .I0(execute_RS2[27]), .I1(_zz_RegFilePlugin_regFile_port1[27]), .S(n3526), .Z(n4220) );
  inv0d0 U6150 ( .I(\RegFilePlugin_regFile[0][26] ), .ZN(n3511) );
  aoi22d1 U6151 ( .A1(n3511), .A2(n3555), .B1(n3510), .B2(n3545), .ZN(n4219)
         );
  mx02d1 U6152 ( .I0(execute_RS1[26]), .I1(_zz_RegFilePlugin_regFile_port0[26]), .S(n3526), .Z(n4218) );
  mx02d1 U6153 ( .I0(execute_RS2[26]), .I1(_zz_RegFilePlugin_regFile_port1[26]), .S(n3516), .Z(n4217) );
  inv0d0 U6154 ( .I(\RegFilePlugin_regFile[0][25] ), .ZN(n3513) );
  aoi22d1 U6155 ( .A1(n3513), .A2(n3555), .B1(n3512), .B2(n3545), .ZN(n4216)
         );
  mx02d1 U6156 ( .I0(execute_RS1[25]), .I1(_zz_RegFilePlugin_regFile_port0[25]), .S(n3516), .Z(n4215) );
  mx02d1 U6157 ( .I0(execute_RS2[25]), .I1(_zz_RegFilePlugin_regFile_port1[25]), .S(n3526), .Z(n4214) );
  inv0d0 U6158 ( .I(\RegFilePlugin_regFile[0][24] ), .ZN(n3514) );
  oai22d1 U6159 ( .A1(n3514), .A2(n3545), .B1(n3341), .B2(n3549), .ZN(n4213)
         );
  mx02d1 U6160 ( .I0(execute_RS1[24]), .I1(_zz_RegFilePlugin_regFile_port0[24]), .S(n3516), .Z(n4212) );
  mx02d1 U6161 ( .I0(execute_RS2[24]), .I1(_zz_RegFilePlugin_regFile_port1[24]), .S(n3526), .Z(n4211) );
  inv0d0 U6162 ( .I(\RegFilePlugin_regFile[0][23] ), .ZN(n3515) );
  aoi22d1 U6163 ( .A1(n3515), .A2(n3555), .B1(n3454), .B2(n3545), .ZN(n4210)
         );
  mx02d1 U6164 ( .I0(execute_RS1[23]), .I1(_zz_RegFilePlugin_regFile_port0[23]), .S(n3539), .Z(n4209) );
  mx02d1 U6165 ( .I0(execute_RS2[23]), .I1(_zz_RegFilePlugin_regFile_port1[23]), .S(n3516), .Z(n4208) );
  inv0d0 U6166 ( .I(\RegFilePlugin_regFile[0][22] ), .ZN(n3518) );
  aoi22d1 U6167 ( .A1(n3518), .A2(n3555), .B1(n3517), .B2(n3556), .ZN(n4207)
         );
  mx02d1 U6168 ( .I0(execute_RS1[22]), .I1(_zz_RegFilePlugin_regFile_port0[22]), .S(n3526), .Z(n4206) );
  mx02d1 U6169 ( .I0(execute_RS2[22]), .I1(_zz_RegFilePlugin_regFile_port1[22]), .S(n3526), .Z(n4205) );
  inv0d0 U6170 ( .I(\RegFilePlugin_regFile[0][21] ), .ZN(n3520) );
  oai22d1 U6171 ( .A1(n3520), .A2(n3556), .B1(n3519), .B2(n3549), .ZN(n4204)
         );
  mx02d1 U6172 ( .I0(execute_RS1[21]), .I1(_zz_RegFilePlugin_regFile_port0[21]), .S(n3526), .Z(n4203) );
  mx02d1 U6173 ( .I0(execute_RS2[21]), .I1(_zz_RegFilePlugin_regFile_port1[21]), .S(n3526), .Z(n4202) );
  inv0d0 U6174 ( .I(\RegFilePlugin_regFile[0][20] ), .ZN(n3522) );
  oai22d1 U6175 ( .A1(n3522), .A2(n3556), .B1(n3521), .B2(n3549), .ZN(n4201)
         );
  mx02d1 U6176 ( .I0(execute_RS1[20]), .I1(_zz_RegFilePlugin_regFile_port0[20]), .S(n3526), .Z(n4200) );
  mx02d1 U6177 ( .I0(execute_RS2[20]), .I1(_zz_RegFilePlugin_regFile_port1[20]), .S(n3526), .Z(n4199) );
  inv0d0 U6178 ( .I(\RegFilePlugin_regFile[0][19] ), .ZN(n3524) );
  oai22d1 U6179 ( .A1(n3524), .A2(n3545), .B1(n3523), .B2(n3555), .ZN(n4198)
         );
  mx02d1 U6180 ( .I0(execute_RS1[19]), .I1(_zz_RegFilePlugin_regFile_port0[19]), .S(n3526), .Z(n4197) );
  mx02d1 U6181 ( .I0(execute_RS2[19]), .I1(_zz_RegFilePlugin_regFile_port1[19]), .S(n3526), .Z(n4196) );
  inv0d0 U6182 ( .I(\RegFilePlugin_regFile[0][18] ), .ZN(n3525) );
  aoi22d1 U6183 ( .A1(n3525), .A2(n3555), .B1(n3456), .B2(n3545), .ZN(n4195)
         );
  mx02d1 U6184 ( .I0(execute_RS1[18]), .I1(_zz_RegFilePlugin_regFile_port0[18]), .S(n3526), .Z(n4194) );
  mx02d1 U6185 ( .I0(execute_RS2[18]), .I1(_zz_RegFilePlugin_regFile_port1[18]), .S(n3539), .Z(n4193) );
  inv0d0 U6186 ( .I(\RegFilePlugin_regFile[0][17] ), .ZN(n3528) );
  aoi22d1 U6187 ( .A1(n3528), .A2(n3549), .B1(n3527), .B2(n3545), .ZN(n4192)
         );
  mx02d1 U6188 ( .I0(execute_RS1[17]), .I1(_zz_RegFilePlugin_regFile_port0[17]), .S(n3548), .Z(n4191) );
  mx02d1 U6189 ( .I0(execute_RS2[17]), .I1(_zz_RegFilePlugin_regFile_port1[17]), .S(n3539), .Z(n4190) );
  inv0d0 U6190 ( .I(\RegFilePlugin_regFile[0][16] ), .ZN(n3530) );
  oai22d1 U6191 ( .A1(n3530), .A2(n3556), .B1(n3529), .B2(n3549), .ZN(n4189)
         );
  mx02d1 U6192 ( .I0(execute_RS1[16]), .I1(_zz_RegFilePlugin_regFile_port0[16]), .S(n3548), .Z(n4188) );
  mx02d1 U6193 ( .I0(execute_RS2[16]), .I1(_zz_RegFilePlugin_regFile_port1[16]), .S(n3548), .Z(n4187) );
  inv0d0 U6194 ( .I(\RegFilePlugin_regFile[0][15] ), .ZN(n3532) );
  aoi22d1 U6195 ( .A1(n3532), .A2(n3555), .B1(n3556), .B2(n3531), .ZN(n4186)
         );
  mx02d1 U6196 ( .I0(execute_RS1[15]), .I1(_zz_RegFilePlugin_regFile_port0[15]), .S(n3539), .Z(n4185) );
  mx02d1 U6197 ( .I0(execute_RS2[15]), .I1(_zz_RegFilePlugin_regFile_port1[15]), .S(n3539), .Z(n4184) );
  inv0d0 U6198 ( .I(\RegFilePlugin_regFile[0][14] ), .ZN(n3533) );
  oai22d1 U6199 ( .A1(n3533), .A2(n3545), .B1(n3459), .B2(n3549), .ZN(n4183)
         );
  mx02d1 U6200 ( .I0(execute_RS1[14]), .I1(_zz_RegFilePlugin_regFile_port0[14]), .S(n3548), .Z(n4182) );
  mx02d1 U6201 ( .I0(execute_RS2[14]), .I1(_zz_RegFilePlugin_regFile_port1[14]), .S(n3539), .Z(n4181) );
  inv0d0 U6202 ( .I(\RegFilePlugin_regFile[0][13] ), .ZN(n3535) );
  aoi22d1 U6203 ( .A1(n3535), .A2(n3555), .B1(n3534), .B2(n3545), .ZN(n4180)
         );
  mx02d1 U6204 ( .I0(execute_RS1[13]), .I1(_zz_RegFilePlugin_regFile_port0[13]), .S(n3539), .Z(n4179) );
  mx02d1 U6205 ( .I0(execute_RS2[13]), .I1(_zz_RegFilePlugin_regFile_port1[13]), .S(n3539), .Z(n4178) );
  inv0d0 U6206 ( .I(\RegFilePlugin_regFile[0][12] ), .ZN(n3536) );
  oai22d1 U6207 ( .A1(n3536), .A2(n3556), .B1(n3460), .B2(n3549), .ZN(n4177)
         );
  mx02d1 U6208 ( .I0(execute_RS1[12]), .I1(_zz_RegFilePlugin_regFile_port0[12]), .S(n3539), .Z(n4176) );
  mx02d1 U6209 ( .I0(execute_RS2[12]), .I1(_zz_RegFilePlugin_regFile_port1[12]), .S(n3539), .Z(n4175) );
  inv0d0 U6210 ( .I(\RegFilePlugin_regFile[0][11] ), .ZN(n3537) );
  oai22d1 U6211 ( .A1(n3537), .A2(n3556), .B1(n3461), .B2(n3549), .ZN(n4174)
         );
  mx02d1 U6212 ( .I0(execute_RS1[11]), .I1(_zz_RegFilePlugin_regFile_port0[11]), .S(n3539), .Z(n4173) );
  mx02d1 U6213 ( .I0(execute_RS2[11]), .I1(_zz_RegFilePlugin_regFile_port1[11]), .S(n3539), .Z(n4172) );
  inv0d0 U6214 ( .I(\RegFilePlugin_regFile[0][10] ), .ZN(n3538) );
  oai22d1 U6215 ( .A1(n3538), .A2(n3545), .B1(n3462), .B2(n3549), .ZN(n4171)
         );
  mx02d1 U6216 ( .I0(execute_RS1[10]), .I1(_zz_RegFilePlugin_regFile_port0[10]), .S(n3539), .Z(n4170) );
  mx02d1 U6217 ( .I0(execute_RS2[10]), .I1(_zz_RegFilePlugin_regFile_port1[10]), .S(n3539), .Z(n4169) );
  inv0d0 U6218 ( .I(\RegFilePlugin_regFile[0][9] ), .ZN(n3540) );
  oai22d1 U6219 ( .A1(n3540), .A2(n3556), .B1(n3463), .B2(n3549), .ZN(n4168)
         );
  mx02d1 U6220 ( .I0(execute_RS1[9]), .I1(_zz_RegFilePlugin_regFile_port0[9]), 
        .S(n3548), .Z(n4167) );
  mx02d1 U6221 ( .I0(execute_RS2[9]), .I1(_zz_RegFilePlugin_regFile_port1[9]), 
        .S(n3548), .Z(n4166) );
  inv0d0 U6222 ( .I(\RegFilePlugin_regFile[0][8] ), .ZN(n3542) );
  oai22d1 U6223 ( .A1(n3542), .A2(n3556), .B1(n3541), .B2(n3549), .ZN(n4165)
         );
  mx02d1 U6224 ( .I0(execute_RS1[8]), .I1(_zz_RegFilePlugin_regFile_port0[8]), 
        .S(n3548), .Z(n4164) );
  mx02d1 U6225 ( .I0(execute_RS2[8]), .I1(_zz_RegFilePlugin_regFile_port1[8]), 
        .S(n3548), .Z(n4163) );
  inv0d0 U6226 ( .I(\RegFilePlugin_regFile[0][7] ), .ZN(n3544) );
  oai22d1 U6227 ( .A1(n3544), .A2(n3556), .B1(n3555), .B2(n3543), .ZN(n4162)
         );
  mx02d1 U6228 ( .I0(execute_RS1[7]), .I1(_zz_RegFilePlugin_regFile_port0[7]), 
        .S(n3548), .Z(n4161) );
  mx02d1 U6229 ( .I0(execute_RS2[7]), .I1(_zz_RegFilePlugin_regFile_port1[7]), 
        .S(n3548), .Z(n4160) );
  inv0d0 U6230 ( .I(\RegFilePlugin_regFile[0][6] ), .ZN(n3546) );
  oai22d1 U6231 ( .A1(n3546), .A2(n3545), .B1(n3555), .B2(n3467), .ZN(n4159)
         );
  mx02d1 U6232 ( .I0(execute_RS1[6]), .I1(_zz_RegFilePlugin_regFile_port0[6]), 
        .S(n3548), .Z(n4158) );
  mx02d1 U6233 ( .I0(execute_RS2[6]), .I1(_zz_RegFilePlugin_regFile_port1[6]), 
        .S(n3548), .Z(n4157) );
  inv0d0 U6234 ( .I(\RegFilePlugin_regFile[0][5] ), .ZN(n3547) );
  oai22d1 U6235 ( .A1(n3547), .A2(n3556), .B1(n3549), .B2(n3468), .ZN(n4156)
         );
  mx02d1 U6236 ( .I0(execute_RS1[5]), .I1(_zz_RegFilePlugin_regFile_port0[5]), 
        .S(n3548), .Z(n4155) );
  mx02d1 U6237 ( .I0(execute_RS2[5]), .I1(_zz_RegFilePlugin_regFile_port1[5]), 
        .S(n3558), .Z(n4154) );
  inv0d0 U6238 ( .I(\RegFilePlugin_regFile[0][4] ), .ZN(n3550) );
  oai22d1 U6239 ( .A1(n3550), .A2(n3556), .B1(n3549), .B2(n3469), .ZN(n4153)
         );
  mx02d1 U6240 ( .I0(execute_RS1[4]), .I1(_zz_RegFilePlugin_regFile_port0[4]), 
        .S(n3558), .Z(n4152) );
  mx02d1 U6241 ( .I0(execute_RS2[4]), .I1(_zz_RegFilePlugin_regFile_port1[4]), 
        .S(n3558), .Z(n4151) );
  inv0d0 U6242 ( .I(\RegFilePlugin_regFile[0][3] ), .ZN(n3552) );
  oai22d1 U6243 ( .A1(n3552), .A2(n3556), .B1(n3555), .B2(n3551), .ZN(n4150)
         );
  mx02d1 U6244 ( .I0(execute_RS1[3]), .I1(_zz_RegFilePlugin_regFile_port0[3]), 
        .S(n3558), .Z(n4149) );
  mx02d1 U6245 ( .I0(execute_RS2[3]), .I1(_zz_RegFilePlugin_regFile_port1[3]), 
        .S(n3558), .Z(n4148) );
  inv0d0 U6246 ( .I(\RegFilePlugin_regFile[0][2] ), .ZN(n3553) );
  oai22d1 U6247 ( .A1(n3553), .A2(n3556), .B1(n3555), .B2(n3472), .ZN(n4147)
         );
  mx02d1 U6248 ( .I0(execute_RS1[2]), .I1(_zz_RegFilePlugin_regFile_port0[2]), 
        .S(n3558), .Z(n4146) );
  mx02d1 U6249 ( .I0(execute_RS2[2]), .I1(_zz_RegFilePlugin_regFile_port1[2]), 
        .S(n3558), .Z(n4145) );
  inv0d0 U6250 ( .I(\RegFilePlugin_regFile[0][1] ), .ZN(n3557) );
  oai22d1 U6251 ( .A1(n3557), .A2(n3556), .B1(n3555), .B2(n3554), .ZN(n4144)
         );
  mx02d1 U6252 ( .I0(execute_RS1[1]), .I1(_zz_RegFilePlugin_regFile_port0[1]), 
        .S(n3558), .Z(n4143) );
  mx02d1 U6253 ( .I0(execute_RS2[1]), .I1(_zz_RegFilePlugin_regFile_port1[1]), 
        .S(n3559), .Z(n4142) );
  nr02d1 U6254 ( .A1(n3561), .A2(n3560), .ZN(n3562) );
  buffd1 U6255 ( .I(n3562), .Z(n3565) );
  aoim22d1 U6256 ( .A1(n3565), .A2(n3573), .B1(CsrPlugin_mtvec_base[0]), .B2(
        n3562), .Z(n4141) );
  buffd1 U6257 ( .I(n3562), .Z(n3564) );
  aoim22d1 U6258 ( .A1(n3565), .A2(n3576), .B1(CsrPlugin_mtvec_base[1]), .B2(
        n3564), .Z(n4140) );
  buffd1 U6259 ( .I(n3562), .Z(n3563) );
  aoim22d1 U6260 ( .A1(n3565), .A2(n3579), .B1(CsrPlugin_mtvec_base[2]), .B2(
        n3563), .Z(n4139) );
  aoim22d1 U6261 ( .A1(n3565), .A2(n3582), .B1(CsrPlugin_mtvec_base[3]), .B2(
        n3564), .Z(n4138) );
  aoim22d1 U6262 ( .A1(n3565), .A2(n3585), .B1(CsrPlugin_mtvec_base[4]), .B2(
        n3564), .Z(n4137) );
  aoim22d1 U6263 ( .A1(n3565), .A2(n3588), .B1(CsrPlugin_mtvec_base[5]), .B2(
        n3563), .Z(n4136) );
  aoim22d1 U6264 ( .A1(n3565), .A2(n3591), .B1(CsrPlugin_mtvec_base[6]), .B2(
        n3563), .Z(n4135) );
  aoim22d1 U6265 ( .A1(n3565), .A2(n3594), .B1(CsrPlugin_mtvec_base[7]), .B2(
        n3563), .Z(n4134) );
  aoim22d1 U6266 ( .A1(n3563), .A2(n3597), .B1(CsrPlugin_mtvec_base[8]), .B2(
        n3563), .Z(n4133) );
  aoim22d1 U6267 ( .A1(n3562), .A2(n3600), .B1(CsrPlugin_mtvec_base[9]), .B2(
        n3563), .Z(n4132) );
  aoim22d1 U6268 ( .A1(n3562), .A2(n3603), .B1(CsrPlugin_mtvec_base[10]), .B2(
        n3563), .Z(n4131) );
  aoim22d1 U6269 ( .A1(n3563), .A2(n3606), .B1(CsrPlugin_mtvec_base[11]), .B2(
        n3563), .Z(n4130) );
  aoim22d1 U6270 ( .A1(n3563), .A2(n3609), .B1(CsrPlugin_mtvec_base[12]), .B2(
        n3563), .Z(n4129) );
  aoim22d1 U6271 ( .A1(n3564), .A2(n3612), .B1(CsrPlugin_mtvec_base[13]), .B2(
        n3563), .Z(n4128) );
  aoim22d1 U6272 ( .A1(n3565), .A2(n3615), .B1(CsrPlugin_mtvec_base[14]), .B2(
        n3563), .Z(n4127) );
  aoim22d1 U6273 ( .A1(n3565), .A2(n3618), .B1(CsrPlugin_mtvec_base[15]), .B2(
        n3562), .Z(n4126) );
  aoim22d1 U6274 ( .A1(n3564), .A2(n3621), .B1(CsrPlugin_mtvec_base[16]), .B2(
        n3563), .Z(n4125) );
  aoim22d1 U6275 ( .A1(n3564), .A2(n3624), .B1(CsrPlugin_mtvec_base[17]), .B2(
        n3562), .Z(n4124) );
  aoim22d1 U6276 ( .A1(n3564), .A2(n3627), .B1(CsrPlugin_mtvec_base[18]), .B2(
        n3562), .Z(n4123) );
  aoim22d1 U6277 ( .A1(n3565), .A2(n3630), .B1(CsrPlugin_mtvec_base[19]), .B2(
        n3564), .Z(n4122) );
  aoim22d1 U6278 ( .A1(n3564), .A2(n3632), .B1(CsrPlugin_mtvec_base[20]), .B2(
        n3562), .Z(n4121) );
  aoim22d1 U6279 ( .A1(n3565), .A2(n3636), .B1(CsrPlugin_mtvec_base[21]), .B2(
        n3562), .Z(n4120) );
  aoim22d1 U6280 ( .A1(n3563), .A2(n3638), .B1(CsrPlugin_mtvec_base[22]), .B2(
        n3562), .Z(n4119) );
  aoim22d1 U6281 ( .A1(n3564), .A2(n3643), .B1(CsrPlugin_mtvec_base[23]), .B2(
        n3564), .Z(n4118) );
  aoim22d1 U6282 ( .A1(n3565), .A2(n3646), .B1(CsrPlugin_mtvec_base[24]), .B2(
        n3562), .Z(n4117) );
  aoim22d1 U6283 ( .A1(n3564), .A2(n3649), .B1(CsrPlugin_mtvec_base[25]), .B2(
        n3564), .Z(n4116) );
  aoim22d1 U6284 ( .A1(n3563), .A2(n3652), .B1(CsrPlugin_mtvec_base[26]), .B2(
        n3564), .Z(n4115) );
  aoim22d1 U6285 ( .A1(n3565), .A2(n3655), .B1(CsrPlugin_mtvec_base[27]), .B2(
        n3564), .Z(n4114) );
  aoim22d1 U6286 ( .A1(n3565), .A2(n3661), .B1(CsrPlugin_mtvec_base[28]), .B2(
        n3564), .Z(n4113) );
  aoim22d1 U6287 ( .A1(n3565), .A2(n3667), .B1(CsrPlugin_mtvec_base[29]), .B2(
        n3564), .Z(n4112) );
  buffd1 U6288 ( .I(n3666), .Z(n3660) );
  buffd1 U6289 ( .I(n3666), .Z(n3642) );
  nd02d1 U6290 ( .A1(n3677), .A2(n3642), .ZN(n3665) );
  buffd1 U6291 ( .I(n3665), .Z(n3659) );
  inv0d0 U6292 ( .I(CsrPlugin_mepc[0]), .ZN(n3567) );
  oai22d1 U6293 ( .A1(n3660), .A2(n3568), .B1(n3659), .B2(n3567), .ZN(n4111)
         );
  oai22d1 U6294 ( .A1(n3660), .A2(n3570), .B1(n3659), .B2(n3569), .ZN(n4110)
         );
  inv0d0 U6295 ( .I(CsrPlugin_mepc[2]), .ZN(n3572) );
  nd02d1 U6296 ( .A1(n3672), .A2(n3642), .ZN(n3656) );
  buffd1 U6297 ( .I(n3656), .Z(n3662) );
  oai222d1 U6298 ( .A1(n3573), .A2(n3642), .B1(n3659), .B2(n3572), .C1(n3662), 
        .C2(n3571), .ZN(n4109) );
  inv0d0 U6299 ( .I(CsrPlugin_mepc[3]), .ZN(n3575) );
  oai222d1 U6300 ( .A1(n3576), .A2(n3642), .B1(n3665), .B2(n3575), .C1(n3662), 
        .C2(n3574), .ZN(n4108) );
  inv0d0 U6301 ( .I(CsrPlugin_mepc[4]), .ZN(n3578) );
  oai222d1 U6302 ( .A1(n3579), .A2(n3642), .B1(n3665), .B2(n3578), .C1(n3662), 
        .C2(n3577), .ZN(n4107) );
  inv0d0 U6303 ( .I(CsrPlugin_mepc[5]), .ZN(n3581) );
  oai222d1 U6304 ( .A1(n3582), .A2(n3642), .B1(n3665), .B2(n3581), .C1(n3580), 
        .C2(n3662), .ZN(n4106) );
  inv0d0 U6305 ( .I(CsrPlugin_mepc[6]), .ZN(n3584) );
  oai222d1 U6306 ( .A1(n3585), .A2(n3642), .B1(n3665), .B2(n3584), .C1(n3583), 
        .C2(n3662), .ZN(n4105) );
  inv0d0 U6307 ( .I(CsrPlugin_mepc[7]), .ZN(n3587) );
  oai222d1 U6308 ( .A1(n3588), .A2(n3660), .B1(n3659), .B2(n3587), .C1(n3662), 
        .C2(n3586), .ZN(n4104) );
  oai222d1 U6309 ( .A1(n3591), .A2(n3660), .B1(n3659), .B2(n3590), .C1(n3589), 
        .C2(n3662), .ZN(n4103) );
  oai222d1 U6310 ( .A1(n3594), .A2(n3660), .B1(n3665), .B2(n3593), .C1(n3592), 
        .C2(n3656), .ZN(n4102) );
  oai222d1 U6311 ( .A1(n3597), .A2(n3660), .B1(n3659), .B2(n3596), .C1(n3595), 
        .C2(n3656), .ZN(n4101) );
  inv0d0 U6312 ( .I(CsrPlugin_mepc[11]), .ZN(n3599) );
  oai222d1 U6313 ( .A1(n3600), .A2(n3660), .B1(n3665), .B2(n3599), .C1(n3662), 
        .C2(n3598), .ZN(n4100) );
  inv0d0 U6314 ( .I(CsrPlugin_mepc[12]), .ZN(n3602) );
  oai222d1 U6315 ( .A1(n3603), .A2(n3660), .B1(n3659), .B2(n3602), .C1(n3662), 
        .C2(n3601), .ZN(n4099) );
  oai222d1 U6316 ( .A1(n3606), .A2(n3666), .B1(n3665), .B2(n3605), .C1(n3604), 
        .C2(n3662), .ZN(n4098) );
  oai222d1 U6317 ( .A1(n3609), .A2(n3642), .B1(n3665), .B2(n3608), .C1(n3607), 
        .C2(n3656), .ZN(n4097) );
  oai222d1 U6318 ( .A1(n3612), .A2(n3660), .B1(n3665), .B2(n3611), .C1(n3610), 
        .C2(n3656), .ZN(n4096) );
  oai222d1 U6319 ( .A1(n3615), .A2(n3666), .B1(n3665), .B2(n3614), .C1(n3613), 
        .C2(n3656), .ZN(n4095) );
  oai222d1 U6320 ( .A1(n3618), .A2(n3666), .B1(n3659), .B2(n3617), .C1(n3662), 
        .C2(n3616), .ZN(n4094) );
  oai222d1 U6321 ( .A1(n3621), .A2(n3666), .B1(n3659), .B2(n3620), .C1(n3619), 
        .C2(n3656), .ZN(n4093) );
  oai222d1 U6322 ( .A1(n3624), .A2(n3660), .B1(n3665), .B2(n3623), .C1(n3622), 
        .C2(n3656), .ZN(n4092) );
  oai222d1 U6323 ( .A1(n3627), .A2(n3666), .B1(n3665), .B2(n3626), .C1(n3625), 
        .C2(n3656), .ZN(n4091) );
  oai222d1 U6324 ( .A1(n3630), .A2(n3642), .B1(n3665), .B2(n3629), .C1(n3628), 
        .C2(n3656), .ZN(n4090) );
  inv0d0 U6325 ( .I(CsrPlugin_mepc[22]), .ZN(n3631) );
  oai222d1 U6326 ( .A1(n3633), .A2(n3662), .B1(n3660), .B2(n3632), .C1(n3631), 
        .C2(n3659), .ZN(n4089) );
  oai222d1 U6327 ( .A1(n3636), .A2(n3666), .B1(n3659), .B2(n3635), .C1(n3634), 
        .C2(n3656), .ZN(n4088) );
  inv0d0 U6328 ( .I(CsrPlugin_mepc[24]), .ZN(n3637) );
  oai222d1 U6329 ( .A1(n3639), .A2(n3656), .B1(n3660), .B2(n3638), .C1(n3637), 
        .C2(n3659), .ZN(n4087) );
  inv0d0 U6330 ( .I(CsrPlugin_mepc[25]), .ZN(n3641) );
  oai222d1 U6331 ( .A1(n3643), .A2(n3642), .B1(n3665), .B2(n3641), .C1(n3640), 
        .C2(n3656), .ZN(n4086) );
  inv0d0 U6332 ( .I(CsrPlugin_mepc[26]), .ZN(n3645) );
  oai222d1 U6333 ( .A1(n3646), .A2(n3660), .B1(n3659), .B2(n3645), .C1(n3644), 
        .C2(n3662), .ZN(n4085) );
  oai222d1 U6334 ( .A1(n3649), .A2(n3660), .B1(n3659), .B2(n3648), .C1(n3647), 
        .C2(n3662), .ZN(n4084) );
  oai222d1 U6335 ( .A1(n3652), .A2(n3660), .B1(n3659), .B2(n3651), .C1(n3650), 
        .C2(n3662), .ZN(n4083) );
  oai222d1 U6336 ( .A1(n3655), .A2(n3660), .B1(n3659), .B2(n3654), .C1(n3653), 
        .C2(n3662), .ZN(n4082) );
  oai222d1 U6337 ( .A1(n3661), .A2(n3660), .B1(n3659), .B2(n3658), .C1(n3657), 
        .C2(n3656), .ZN(n4081) );
  inv0d0 U6338 ( .I(CsrPlugin_mepc[31]), .ZN(n3664) );
  oai222d1 U6339 ( .A1(n3667), .A2(n3666), .B1(n3665), .B2(n3664), .C1(n3663), 
        .C2(n3662), .ZN(n4080) );
  oaim21d1 U6340 ( .B1(n3669), .B2(\CsrPlugin_interrupt_code[3] ), .A(n3668), 
        .ZN(n4078) );
  aoim22d1 U6341 ( .A1(n3671), .A2(n3670), .B1(
        CsrPlugin_mcause_exceptionCode[0]), .B2(n3672), .Z(n4077) );
  oai22d1 U6342 ( .A1(n3673), .A2(
        CsrPlugin_exceptionPortCtrl_exceptionContext_code[1]), .B1(
        CsrPlugin_mcause_exceptionCode[1]), .B2(n3672), .ZN(n3674) );
  inv0d0 U6343 ( .I(n3674), .ZN(n4076) );
  aor222d1 U6344 ( .A1(CsrPlugin_mcause_exceptionCode[3]), .A2(n3677), .B1(
        CsrPlugin_exceptionPortCtrl_exceptionContext_code[3]), .B2(n3676), 
        .C1(n3675), .C2(\CsrPlugin_interrupt_code[3] ), .Z(n4074) );
  oai22d1 U6345 ( .A1(n3679), .A2(execute_LightShifterPlugin_amplitudeReg[0]), 
        .B1(n3678), .B2(execute_LightShifterPlugin_isActive), .ZN(n3682) );
  inv0d0 U6346 ( .I(n3682), .ZN(n3699) );
  aoim22d1 U6347 ( .A1(n3697), .A2(n3699), .B1(
        execute_LightShifterPlugin_amplitudeReg[0]), .B2(n3697), .Z(n4073) );
  aoi22d1 U6348 ( .A1(n3680), .A2(n3682), .B1(n3699), .B2(n3686), .ZN(n3681)
         );
  aoim22d1 U6349 ( .A1(n3697), .A2(n3681), .B1(
        execute_LightShifterPlugin_amplitudeReg[1]), .B2(n3697), .Z(n4072) );
  nd02d0 U6350 ( .A1(n3683), .A2(n3682), .ZN(n3691) );
  inv0d0 U6351 ( .I(n3691), .ZN(n3684) );
  oan211d1 U6352 ( .C1(n3686), .C2(n3699), .B(n3685), .A(n3684), .ZN(n3689) );
  aoi22d1 U6353 ( .A1(n3697), .A2(n3689), .B1(n3688), .B2(n3687), .ZN(n4071)
         );
  inv0d0 U6354 ( .I(n3690), .ZN(n3692) );
  oai21d1 U6355 ( .B1(n3692), .B2(n3691), .A(n3697), .ZN(n3696) );
  aoi21d1 U6356 ( .B1(n3692), .B2(n3691), .A(n3696), .ZN(n3693) );
  aoim21d1 U6357 ( .B1(execute_LightShifterPlugin_amplitudeReg[3]), .B2(n3697), 
        .A(n3693), .ZN(n4070) );
  inv0d0 U6358 ( .I(n3694), .ZN(n3700) );
  inv0d0 U6359 ( .I(execute_LightShifterPlugin_amplitudeReg[4]), .ZN(n3698) );
  oai222d1 U6360 ( .A1(n3700), .A2(n3699), .B1(n3698), .B2(n3697), .C1(n3696), 
        .C2(n3695), .ZN(n4069) );
  aon211d1 U6361 ( .C1(debug_bus_cmd_payload_data[16]), .C2(n3703), .B(
        DebugPlugin_resetIt), .A(n3701), .ZN(n3702) );
  aoi21d1 U6362 ( .B1(debug_bus_cmd_payload_data[24]), .B2(n3703), .A(n3702), 
        .ZN(n4068) );
  nr02d0 U6363 ( .A1(n3705), .A2(n3706), .ZN(n3704) );
  nd02d0 U6364 ( .A1(n3710), .A2(n3704), .ZN(n3707) );
  nr02d1 U6365 ( .A1(n7005), .A2(n3707), .ZN(n6772) );
  buffd1 U6366 ( .I(n6772), .Z(n7096) );
  nd02d0 U6367 ( .A1(n3710), .A2(n3722), .ZN(n3720) );
  nr02d1 U6368 ( .A1(n7005), .A2(n3720), .ZN(n6465) );
  buffd1 U6369 ( .I(n6465), .Z(n6754) );
  aoi22d1 U6370 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][31] ), 
        .B1(n6754), .B2(\IBusCachedPlugin_cache/banks_0[3][31] ), .ZN(n3716)
         );
  inv0d0 U6371 ( .I(n3710), .ZN(n3721) );
  nd02d0 U6372 ( .A1(n3704), .A2(n3721), .ZN(n3725) );
  nr02d1 U6373 ( .A1(n7005), .A2(n3725), .ZN(n6628) );
  buffd1 U6374 ( .I(n6628), .Z(n6599) );
  inv0d0 U6375 ( .I(n3705), .ZN(n3708) );
  nr02d0 U6376 ( .A1(n3708), .A2(n3706), .ZN(n3717) );
  nd02d0 U6377 ( .A1(n3710), .A2(n3717), .ZN(n3718) );
  buffd1 U6378 ( .I(n6460), .Z(n6789) );
  aoi22d1 U6379 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][31] ), 
        .B1(n6789), .B2(\IBusCachedPlugin_cache/banks_0[0][31] ), .ZN(n3715)
         );
  nr02d1 U6380 ( .A1(n7006), .A2(n3707), .ZN(n6438) );
  buffd1 U6381 ( .I(n6438), .Z(n7097) );
  nd02d0 U6382 ( .A1(n3710), .A2(n3711), .ZN(n3719) );
  nr02d1 U6383 ( .A1(n7005), .A2(n3719), .ZN(n6767) );
  buffd1 U6384 ( .I(n6767), .Z(n6783) );
  aoi22d1 U6385 ( .A1(n7097), .A2(\IBusCachedPlugin_cache/banks_0[10][31] ), 
        .B1(n6783), .B2(\IBusCachedPlugin_cache/banks_0[1][31] ), .ZN(n3714)
         );
  nd02d0 U6386 ( .A1(n3711), .A2(n3721), .ZN(n3712) );
  nr02d1 U6387 ( .A1(n7005), .A2(n3712), .ZN(n6637) );
  buffd1 U6388 ( .I(n6637), .Z(n6791) );
  aoi22d1 U6389 ( .A1(n6791), .A2(\IBusCachedPlugin_cache/banks_0[5][31] ), 
        .B1(n6672), .B2(\IBusCachedPlugin_cache/banks_0[13][31] ), .ZN(n3713)
         );
  nd02d0 U6390 ( .A1(n3717), .A2(n3721), .ZN(n3724) );
  nr02d1 U6391 ( .A1(n7005), .A2(n3724), .ZN(n6554) );
  buffd1 U6392 ( .I(n6554), .Z(n7102) );
  buffd1 U6393 ( .I(n6528), .Z(n7095) );
  aoi22d1 U6394 ( .A1(n7102), .A2(\IBusCachedPlugin_cache/banks_0[4][31] ), 
        .B1(n7095), .B2(\IBusCachedPlugin_cache/banks_0[8][31] ), .ZN(n3729)
         );
  nr02d1 U6395 ( .A1(n7006), .A2(n3720), .ZN(n6652) );
  buffd1 U6396 ( .I(n6652), .Z(n6784) );
  aoi22d1 U6397 ( .A1(n6651), .A2(\IBusCachedPlugin_cache/banks_0[9][31] ), 
        .B1(n6784), .B2(\IBusCachedPlugin_cache/banks_0[11][31] ), .ZN(n3728)
         );
  nd02d0 U6398 ( .A1(n3722), .A2(n3721), .ZN(n3723) );
  nr02d1 U6399 ( .A1(n7005), .A2(n3723), .ZN(n6247) );
  buffd1 U6400 ( .I(n6247), .Z(n6723) );
  nr02d1 U6401 ( .A1(n7006), .A2(n3723), .ZN(n6671) );
  buffd1 U6402 ( .I(n6671), .Z(n6729) );
  aoi22d1 U6403 ( .A1(n6723), .A2(\IBusCachedPlugin_cache/banks_0[7][31] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][31] ), .ZN(n3727)
         );
  nr02d1 U6404 ( .A1(n7006), .A2(n3724), .ZN(n6475) );
  buffd1 U6405 ( .I(n6475), .Z(n6790) );
  nr02d1 U6406 ( .A1(n7006), .A2(n3725), .ZN(n6537) );
  buffd1 U6407 ( .I(n6537), .Z(n6696) );
  aoi22d1 U6408 ( .A1(n6790), .A2(\IBusCachedPlugin_cache/banks_0[12][31] ), 
        .B1(n6696), .B2(\IBusCachedPlugin_cache/banks_0[14][31] ), .ZN(n3726)
         );
  inv0d1 U6409 ( .I(n6936), .ZN(n7107) );
  oai21d1 U6410 ( .B1(n3731), .B2(n3730), .A(n7107), .ZN(n3732) );
  oai21d1 U6411 ( .B1(n7007), .B2(n3733), .A(n3732), .ZN(n4067) );
  nr04d0 U6412 ( .A1(n3737), .A2(n3736), .A3(n3735), .A4(n3734), .ZN(n3776) );
  nr04d0 U6413 ( .A1(n3741), .A2(n3740), .A3(n3739), .A4(n3738), .ZN(n3775) );
  nr04d0 U6414 ( .A1(n3745), .A2(n3744), .A3(n3743), .A4(n3742), .ZN(n3747) );
  oai211d1 U6415 ( .C1(n3749), .C2(n3748), .A(n3747), .B(n3746), .ZN(n3771) );
  nr04d0 U6416 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3769) );
  nr04d0 U6417 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3768) );
  nr04d0 U6418 ( .A1(n3761), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n3767) );
  nr04d0 U6419 ( .A1(n3765), .A2(n3764), .A3(n3763), .A4(n3762), .ZN(n3766) );
  oai21d1 U6420 ( .B1(n3778), .B2(n6681), .A(n6666), .ZN(n3777) );
  aon211d1 U6421 ( .C1(n3778), .C2(n6681), .B(n3777), .A(n6650), .ZN(n3781) );
  aoi21d1 U6422 ( .B1(n3782), .B2(n6681), .A(n6650), .ZN(n3779) );
  oan211d1 U6423 ( .C1(n3782), .C2(n6681), .B(n3779), .A(n6268), .ZN(n3780) );
  aon211d1 U6424 ( .C1(n3782), .C2(
        _zz__zz_execute_BranchPlugin_branch_src2[12]), .B(n3781), .A(n3780), 
        .ZN(n3784) );
  inv0d1 U6425 ( .I(n7113), .ZN(n7120) );
  nd02d0 U6426 ( .A1(n7120), .A2(memory_BRANCH_DO), .ZN(n3783) );
  aon211d1 U6427 ( .C1(n3784), .C2(n6302), .B(n6740), .A(n3783), .ZN(n4066) );
  inv0d0 U6428 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[26] ), .ZN(
        n7015) );
  oai22d1 U6429 ( .A1(n6869), .A2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[13] ), .B1(n7015), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[30]), .ZN(n3785) );
  aoi221d1 U6430 ( .B1(n6869), .B2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[13] ), .C1(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[30]), .C2(n7015), .A(
        n3785), .ZN(n3815) );
  inv0d0 U6431 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[20] ), .ZN(
        n7033) );
  oai22d1 U6432 ( .A1(n6892), .A2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[9] ), .B1(n7033), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[24]), .ZN(n3786) );
  aoi221d1 U6433 ( .B1(n6892), .B2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[9] ), .C1(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[24]), .C2(n7033), .A(
        n3786), .ZN(n3814) );
  inv0d0 U6434 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[22] ), .ZN(
        n7027) );
  aoi22d1 U6435 ( .A1(IBusCachedPlugin_iBusRsp_stages_1_input_payload[26]), 
        .A2(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[22] ), .B1(n7027), 
        .B2(n6823), .ZN(n3790) );
  inv0d0 U6436 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[2] ), .ZN(
        n7091) );
  aoi22d1 U6437 ( .A1(IBusCachedPlugin_iBusRsp_stages_1_input_payload[6]), 
        .A2(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[2] ), .B1(n7091), 
        .B2(n6938), .ZN(n3789) );
  inv0d0 U6438 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[7] ), .ZN(
        n7072) );
  aoi22d1 U6439 ( .A1(IBusCachedPlugin_iBusRsp_stages_1_input_payload[11]), 
        .A2(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[7] ), .B1(n7072), 
        .B2(n6899), .ZN(n3788) );
  inv0d0 U6440 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[14] ), .ZN(
        n7051) );
  aoi22d1 U6441 ( .A1(IBusCachedPlugin_iBusRsp_stages_1_input_payload[18]), 
        .A2(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[14] ), .B1(n7051), 
        .B2(n6864), .ZN(n3787) );
  nr04d0 U6442 ( .A1(n3790), .A2(n3789), .A3(n3788), .A4(n3787), .ZN(n3813) );
  inv0d0 U6443 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[17] ), .ZN(
        n7042) );
  aoi22d1 U6444 ( .A1(IBusCachedPlugin_iBusRsp_stages_1_input_payload[21]), 
        .A2(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[17] ), .B1(n7042), 
        .B2(n6848), .ZN(n3811) );
  inv0d0 U6445 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[8] ), .ZN(
        n7069) );
  aoi22d1 U6446 ( .A1(IBusCachedPlugin_iBusRsp_stages_1_input_payload[12]), 
        .A2(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[8] ), .B1(n7069), 
        .B2(n3820), .ZN(n3810) );
  inv0d0 U6447 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[18] ), .ZN(
        n7039) );
  oai22d1 U6448 ( .A1(n6853), .A2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[16] ), .B1(n7039), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[22]), .ZN(n3791) );
  aoi221d1 U6449 ( .B1(n6853), .B2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[16] ), .C1(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[22]), .C2(n7039), .A(
        n3791), .ZN(n3798) );
  inv0d0 U6450 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[10] ), .ZN(
        n7063) );
  oai22d1 U6451 ( .A1(n6925), .A2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[3] ), .B1(n7063), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[14]), .ZN(n3792) );
  aoi221d1 U6452 ( .B1(n6925), .B2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[3] ), .C1(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[14]), .C2(n7063), .A(
        n3792), .ZN(n3797) );
  inv0d0 U6453 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[25] ), .ZN(
        n7018) );
  oai22d1 U6454 ( .A1(n6828), .A2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[21] ), .B1(n7018), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[29]), .ZN(n3793) );
  aoi221d1 U6455 ( .B1(n6828), .B2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[21] ), .C1(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[29]), .C2(n7018), .A(
        n3793), .ZN(n3796) );
  inv0d0 U6456 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[23] ), .ZN(
        n7024) );
  oai22d1 U6457 ( .A1(n6904), .A2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[6] ), .B1(n7024), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[27]), .ZN(n3794) );
  aoi221d1 U6458 ( .B1(n6904), .B2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[6] ), .C1(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[27]), .C2(n7024), .A(
        n3794), .ZN(n3795) );
  inv0d0 U6459 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[19] ), .ZN(
        n7036) );
  oai22d1 U6460 ( .A1(n6874), .A2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[12] ), .B1(n7036), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[23]), .ZN(n3799) );
  aoi221d1 U6461 ( .B1(n6874), .B2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[12] ), .C1(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[23]), .C2(n7036), .A(
        n3799), .ZN(n3807) );
  inv0d0 U6462 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[5] ), .ZN(
        n7079) );
  oai22d1 U6463 ( .A1(n6915), .A2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[4] ), .B1(n7079), .B2(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[9]), .ZN(n3800) );
  aoi221d1 U6464 ( .B1(n6915), .B2(
        \IBusCachedPlugin_cache/_zz_ways_0_tags_port1[4] ), .C1(
        IBusCachedPlugin_iBusRsp_stages_1_input_payload[9]), .C2(n7079), .A(
        n3800), .ZN(n3806) );
  inv0d0 U6465 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[27] ), .ZN(
        n7012) );
  aoi22d1 U6466 ( .A1(IBusCachedPlugin_iBusRsp_stages_1_input_payload[31]), 
        .A2(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[27] ), .B1(n7012), 
        .B2(n3824), .ZN(n3804) );
  inv0d0 U6467 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[15] ), .ZN(
        n7048) );
  aoi22d1 U6468 ( .A1(IBusCachedPlugin_iBusRsp_stages_1_input_payload[19]), 
        .A2(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[15] ), .B1(n7048), 
        .B2(n6858), .ZN(n3803) );
  inv0d0 U6469 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[24] ), .ZN(
        n7021) );
  aoi22d1 U6470 ( .A1(IBusCachedPlugin_iBusRsp_stages_1_input_payload[28]), 
        .A2(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[24] ), .B1(n7021), 
        .B2(n6813), .ZN(n3802) );
  inv0d0 U6471 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[11] ), .ZN(
        n7060) );
  aoi22d1 U6472 ( .A1(IBusCachedPlugin_iBusRsp_stages_1_input_payload[15]), 
        .A2(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[11] ), .B1(n7060), 
        .B2(n6881), .ZN(n3801) );
  nr04d0 U6473 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3805) );
  nr04d0 U6474 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3812) );
  oai22d1 U6475 ( .A1(n3818), .A2(n3817), .B1(n6862), .B2(n3816), .ZN(n4065)
         );
  aoi22d1 U6476 ( .A1(n7085), .A2(n3820), .B1(n3819), .B2(n6862), .ZN(n4064)
         );
  aoi22d1 U6477 ( .A1(n6939), .A2(n3822), .B1(n3821), .B2(n6862), .ZN(n4063)
         );
  aoi22d1 U6478 ( .A1(n6939), .A2(n3824), .B1(n3823), .B2(n6862), .ZN(n4062)
         );
  aoi22d1 U6479 ( .A1(n7120), .A2(n3825), .B1(n6299), .B2(n6996), .ZN(n4060)
         );
  aoi22d1 U6480 ( .A1(n6789), .A2(\IBusCachedPlugin_cache/banks_0[0][0] ), 
        .B1(n6247), .B2(\IBusCachedPlugin_cache/banks_0[7][0] ), .ZN(n3829) );
  aoi22d1 U6481 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][0] ), 
        .B1(n6784), .B2(\IBusCachedPlugin_cache/banks_0[11][0] ), .ZN(n3828)
         );
  aoi22d1 U6482 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][0] ), 
        .B1(n6754), .B2(\IBusCachedPlugin_cache/banks_0[3][0] ), .ZN(n3827) );
  aoi22d1 U6483 ( .A1(n6696), .A2(\IBusCachedPlugin_cache/banks_0[14][0] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][0] ), .ZN(n3826)
         );
  aoi22d1 U6484 ( .A1(n7097), .A2(\IBusCachedPlugin_cache/banks_0[10][0] ), 
        .B1(n6790), .B2(\IBusCachedPlugin_cache/banks_0[12][0] ), .ZN(n4061)
         );
  buffd1 U6485 ( .I(n6528), .Z(n6728) );
  aoi22d1 U6486 ( .A1(n6651), .A2(\IBusCachedPlugin_cache/banks_0[9][0] ), 
        .B1(n6728), .B2(\IBusCachedPlugin_cache/banks_0[8][0] ), .ZN(n4026) );
  aoi22d1 U6487 ( .A1(n6791), .A2(\IBusCachedPlugin_cache/banks_0[5][0] ), 
        .B1(n7102), .B2(\IBusCachedPlugin_cache/banks_0[4][0] ), .ZN(n4022) );
  aoi22d1 U6488 ( .A1(n6772), .A2(\IBusCachedPlugin_cache/banks_0[2][0] ), 
        .B1(n6783), .B2(\IBusCachedPlugin_cache/banks_0[1][0] ), .ZN(n3830) );
  oai21d1 U6489 ( .B1(n5319), .B2(n4079), .A(n7107), .ZN(n5320) );
  oai21d1 U6490 ( .B1(n7007), .B2(n5321), .A(n5320), .ZN(n4059) );
  aoi22d1 U6491 ( .A1(n6475), .A2(\IBusCachedPlugin_cache/banks_0[12][2] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][2] ), .ZN(n6122)
         );
  aoi22d1 U6492 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][2] ), 
        .B1(n6754), .B2(\IBusCachedPlugin_cache/banks_0[3][2] ), .ZN(n6121) );
  aoi22d1 U6493 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][2] ), 
        .B1(n6783), .B2(\IBusCachedPlugin_cache/banks_0[1][2] ), .ZN(n5323) );
  aoi22d1 U6494 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][2] ), 
        .B1(n7095), .B2(\IBusCachedPlugin_cache/banks_0[8][2] ), .ZN(n5322) );
  aoi22d1 U6495 ( .A1(n6651), .A2(\IBusCachedPlugin_cache/banks_0[9][2] ), 
        .B1(n6784), .B2(\IBusCachedPlugin_cache/banks_0[11][2] ), .ZN(n6251)
         );
  aoi22d1 U6496 ( .A1(n6696), .A2(\IBusCachedPlugin_cache/banks_0[14][2] ), 
        .B1(n6247), .B2(\IBusCachedPlugin_cache/banks_0[7][2] ), .ZN(n6250) );
  aoi22d1 U6497 ( .A1(n6791), .A2(\IBusCachedPlugin_cache/banks_0[5][2] ), 
        .B1(n7097), .B2(\IBusCachedPlugin_cache/banks_0[10][2] ), .ZN(n6249)
         );
  aoi22d1 U6498 ( .A1(n6789), .A2(\IBusCachedPlugin_cache/banks_0[0][2] ), 
        .B1(n6554), .B2(\IBusCachedPlugin_cache/banks_0[4][2] ), .ZN(n6248) );
  oai21d1 U6499 ( .B1(n6253), .B2(n6252), .A(n7107), .ZN(n6254) );
  oai21d1 U6500 ( .B1(n7007), .B2(n6255), .A(n6254), .ZN(n4058) );
  an02d1 U6501 ( .A1(execute_BRANCH_CTRL[1]), .A2(execute_BRANCH_CTRL[0]), .Z(
        n6297) );
  buffd1 U6502 ( .I(n6297), .Z(n6301) );
  aoi22d1 U6503 ( .A1(n6301), .A2(n6256), .B1(n6416), .B2(n6290), .ZN(n6310)
         );
  aoi22d1 U6504 ( .A1(n6301), .A2(n6257), .B1(n6418), .B2(n6305), .ZN(n6313)
         );
  aoi22d1 U6505 ( .A1(n6301), .A2(n6258), .B1(n6809), .B2(n6305), .ZN(n6316)
         );
  aoi22d1 U6506 ( .A1(n6301), .A2(n6259), .B1(n6814), .B2(n6290), .ZN(n6319)
         );
  aoi22d1 U6507 ( .A1(n6301), .A2(n6260), .B1(n6819), .B2(n6290), .ZN(n6322)
         );
  aoi22d1 U6508 ( .A1(n6297), .A2(n6261), .B1(n6824), .B2(n6290), .ZN(n6325)
         );
  aoi22d1 U6509 ( .A1(n6301), .A2(n6262), .B1(n6829), .B2(n6290), .ZN(n6328)
         );
  aoi22d1 U6510 ( .A1(n6297), .A2(n6263), .B1(n6834), .B2(n6290), .ZN(n6331)
         );
  aoi22d1 U6511 ( .A1(n6297), .A2(n6264), .B1(n6839), .B2(n6290), .ZN(n6334)
         );
  aoi22d1 U6512 ( .A1(n6297), .A2(n6265), .B1(n6844), .B2(n6290), .ZN(n6337)
         );
  aoi22d1 U6513 ( .A1(n6297), .A2(n6266), .B1(n6849), .B2(n6290), .ZN(n6340)
         );
  aoi22d1 U6514 ( .A1(n6297), .A2(n6267), .B1(n6854), .B2(n6290), .ZN(n6344)
         );
  nd02d1 U6515 ( .A1(execute_BRANCH_CTRL[1]), .A2(n6268), .ZN(n6283) );
  nd02d0 U6516 ( .A1(n6343), .A2(n6283), .ZN(n6281) );
  oai21d1 U6517 ( .B1(n6283), .B2(n6269), .A(n6281), .ZN(n6348) );
  aoi22d1 U6518 ( .A1(n6297), .A2(n6270), .B1(n6859), .B2(n6290), .ZN(n6347)
         );
  oai21d1 U6519 ( .B1(n6283), .B2(n6271), .A(n6281), .ZN(n6352) );
  aoi22d1 U6520 ( .A1(n6301), .A2(n6272), .B1(n6865), .B2(n6290), .ZN(n6351)
         );
  oai21d1 U6521 ( .B1(n6283), .B2(n6273), .A(n6281), .ZN(n6356) );
  aoi22d1 U6522 ( .A1(n6301), .A2(n6274), .B1(n6870), .B2(n6290), .ZN(n6355)
         );
  oai21d1 U6523 ( .B1(n6283), .B2(n6275), .A(n6281), .ZN(n6360) );
  aoi22d1 U6524 ( .A1(n6301), .A2(n6276), .B1(n6875), .B2(n6290), .ZN(n6359)
         );
  oai21d1 U6525 ( .B1(n6283), .B2(n6277), .A(n6281), .ZN(n6364) );
  aoi22d1 U6526 ( .A1(n6301), .A2(n6278), .B1(n6882), .B2(n6290), .ZN(n6363)
         );
  oai21d1 U6527 ( .B1(n6283), .B2(n6650), .A(n6281), .ZN(n6368) );
  aoi22d1 U6528 ( .A1(n6301), .A2(n6279), .B1(n6887), .B2(n6290), .ZN(n6367)
         );
  oai21d1 U6529 ( .B1(n6283), .B2(n6919), .A(n6281), .ZN(n6372) );
  aoi22d1 U6530 ( .A1(n6301), .A2(n6280), .B1(n6894), .B2(n6290), .ZN(n6371)
         );
  oai21d1 U6531 ( .B1(n6283), .B2(n6681), .A(n6281), .ZN(n6376) );
  aoi22d1 U6532 ( .A1(n6301), .A2(n6282), .B1(n7118), .B2(n6290), .ZN(n6375)
         );
  oai222d1 U6533 ( .A1(n6290), .A2(n6284), .B1(n6753), .B2(
        execute_BRANCH_CTRL[1]), .C1(n6307), .C2(n6283), .ZN(n6380) );
  aoi22d1 U6534 ( .A1(n6301), .A2(n6285), .B1(n6900), .B2(n6290), .ZN(n6379)
         );
  aoi22d1 U6535 ( .A1(n6297), .A2(n6286), .B1(n6905), .B2(n6290), .ZN(n6383)
         );
  aoi22d1 U6536 ( .A1(n6297), .A2(n6287), .B1(n6911), .B2(n6290), .ZN(n6386)
         );
  aoi22d1 U6537 ( .A1(n6297), .A2(n6288), .B1(n6916), .B2(n6290), .ZN(n6389)
         );
  aoi22d1 U6538 ( .A1(n6297), .A2(n6289), .B1(n6927), .B2(n6290), .ZN(n6392)
         );
  aoi22d1 U6539 ( .A1(n6297), .A2(n6291), .B1(n6940), .B2(n6290), .ZN(n6395)
         );
  inv0d0 U6540 ( .I(n6301), .ZN(n6305) );
  aoi22d1 U6541 ( .A1(n6297), .A2(n6292), .B1(n7002), .B2(n6305), .ZN(n6398)
         );
  aoi22d1 U6542 ( .A1(execute_BRANCH_CTRL[1]), .A2(n6293), .B1(n6694), .B2(
        n6302), .ZN(n6402) );
  aoi22d1 U6543 ( .A1(n6297), .A2(n6294), .B1(n7114), .B2(n6305), .ZN(n6401)
         );
  aoi22d1 U6544 ( .A1(execute_BRANCH_CTRL[1]), .A2(n6295), .B1(n6709), .B2(
        n6302), .ZN(n6406) );
  aoi22d1 U6545 ( .A1(n6297), .A2(n6296), .B1(n6420), .B2(n6305), .ZN(n6405)
         );
  aoi22d1 U6546 ( .A1(execute_BRANCH_CTRL[1]), .A2(n6298), .B1(n6722), .B2(
        n6302), .ZN(n6410) );
  aoi22d1 U6547 ( .A1(n6301), .A2(n6300), .B1(n6299), .B2(n6305), .ZN(n6409)
         );
  aoi22d1 U6548 ( .A1(execute_BRANCH_CTRL[1]), .A2(n6303), .B1(n6738), .B2(
        n6302), .ZN(n6414) );
  nr02d0 U6549 ( .A1(n6304), .A2(n6305), .ZN(n6413) );
  an02d0 U6550 ( .A1(n6308), .A2(_zz__zz_execute_BranchPlugin_branch_src2[10]), 
        .Z(n6412) );
  xr03d1 U6551 ( .A1(n6310), .A2(n6343), .A3(n6309), .Z(n6311) );
  inv0d0 U6552 ( .I(n6926), .ZN(n6942) );
  mx02d1 U6553 ( .I0(n6311), .I1(memory_BRANCH_CALC[31]), .S(n6942), .Z(n4057)
         );
  mx02d1 U6554 ( .I0(n6314), .I1(memory_BRANCH_CALC[30]), .S(n6889), .Z(n4056)
         );
  inv0d0 U6555 ( .I(n6926), .ZN(n7004) );
  mx02d1 U6556 ( .I0(n6317), .I1(memory_BRANCH_CALC[29]), .S(n7004), .Z(n4055)
         );
  mx02d1 U6557 ( .I0(n6320), .I1(memory_BRANCH_CALC[28]), .S(n6942), .Z(n4054)
         );
  mx02d1 U6558 ( .I0(n6323), .I1(memory_BRANCH_CALC[27]), .S(n7004), .Z(n4053)
         );
  mx02d1 U6559 ( .I0(n6326), .I1(memory_BRANCH_CALC[26]), .S(n7116), .Z(n4052)
         );
  mx02d1 U6560 ( .I0(n6329), .I1(memory_BRANCH_CALC[25]), .S(n6942), .Z(n4051)
         );
  mx02d1 U6561 ( .I0(n6332), .I1(memory_BRANCH_CALC[24]), .S(n7116), .Z(n4050)
         );
  mx02d1 U6562 ( .I0(n6335), .I1(memory_BRANCH_CALC[23]), .S(n7116), .Z(n4049)
         );
  mx02d1 U6563 ( .I0(n6338), .I1(memory_BRANCH_CALC[22]), .S(n6942), .Z(n4048)
         );
  mx02d1 U6564 ( .I0(n6341), .I1(memory_BRANCH_CALC[21]), .S(n6889), .Z(n4047)
         );
  mx02d1 U6565 ( .I0(n6345), .I1(memory_BRANCH_CALC[20]), .S(n7116), .Z(n4046)
         );
  mx02d1 U6566 ( .I0(n6349), .I1(memory_BRANCH_CALC[19]), .S(n7116), .Z(n4045)
         );
  mx02d1 U6567 ( .I0(n6353), .I1(memory_BRANCH_CALC[18]), .S(n7116), .Z(n4044)
         );
  mx02d1 U6568 ( .I0(n6357), .I1(memory_BRANCH_CALC[17]), .S(n7004), .Z(n4043)
         );
  mx02d1 U6569 ( .I0(n6361), .I1(memory_BRANCH_CALC[16]), .S(n6942), .Z(n4042)
         );
  mx02d1 U6570 ( .I0(n6365), .I1(memory_BRANCH_CALC[15]), .S(n7004), .Z(n4041)
         );
  mx02d1 U6571 ( .I0(n6369), .I1(memory_BRANCH_CALC[14]), .S(n6889), .Z(n4040)
         );
  mx02d1 U6572 ( .I0(n6373), .I1(memory_BRANCH_CALC[13]), .S(n7004), .Z(n4039)
         );
  mx02d1 U6573 ( .I0(n6377), .I1(memory_BRANCH_CALC[12]), .S(n7116), .Z(n4038)
         );
  mx02d1 U6574 ( .I0(n6381), .I1(memory_BRANCH_CALC[11]), .S(n7004), .Z(n4037)
         );
  mx02d1 U6575 ( .I0(n6384), .I1(memory_BRANCH_CALC[10]), .S(n7116), .Z(n4036)
         );
  mx02d1 U6576 ( .I0(n6387), .I1(memory_BRANCH_CALC[9]), .S(n7120), .Z(n4035)
         );
  mx02d1 U6577 ( .I0(n6390), .I1(memory_BRANCH_CALC[8]), .S(n7120), .Z(n4034)
         );
  mx02d1 U6578 ( .I0(n6393), .I1(memory_BRANCH_CALC[7]), .S(n7120), .Z(n4033)
         );
  mx02d1 U6579 ( .I0(n6396), .I1(memory_BRANCH_CALC[6]), .S(n6942), .Z(n4032)
         );
  mx02d1 U6580 ( .I0(n6399), .I1(memory_BRANCH_CALC[5]), .S(n7116), .Z(n4031)
         );
  mx02d1 U6581 ( .I0(n6403), .I1(memory_BRANCH_CALC[4]), .S(n7116), .Z(n4030)
         );
  mx02d1 U6582 ( .I0(n6407), .I1(memory_BRANCH_CALC[3]), .S(n7116), .Z(n4029)
         );
  mx02d1 U6583 ( .I0(n6411), .I1(memory_BRANCH_CALC[2]), .S(n6942), .Z(n4028)
         );
  mx02d1 U6584 ( .I0(n6415), .I1(memory_BRANCH_CALC[1]), .S(n7116), .Z(n4027)
         );
  aoi22d1 U6585 ( .A1(n7120), .A2(n6417), .B1(n6416), .B2(n6997), .ZN(n4025)
         );
  aoi22d1 U6586 ( .A1(n6740), .A2(n6419), .B1(n6418), .B2(n7117), .ZN(n4024)
         );
  aoi22d1 U6587 ( .A1(n6740), .A2(n6421), .B1(n6420), .B2(n6997), .ZN(n4023)
         );
  inv0d1 U6588 ( .I(n6936), .ZN(n7112) );
  aoi22d1 U6589 ( .A1(n6438), .A2(\IBusCachedPlugin_cache/banks_0[10][3] ), 
        .B1(n6475), .B2(\IBusCachedPlugin_cache/banks_0[12][3] ), .ZN(n6425)
         );
  aoi22d1 U6590 ( .A1(n6460), .A2(\IBusCachedPlugin_cache/banks_0[0][3] ), 
        .B1(n6784), .B2(\IBusCachedPlugin_cache/banks_0[11][3] ), .ZN(n6424)
         );
  aoi22d1 U6591 ( .A1(n6651), .A2(\IBusCachedPlugin_cache/banks_0[9][3] ), 
        .B1(n7095), .B2(\IBusCachedPlugin_cache/banks_0[8][3] ), .ZN(n6423) );
  aoi22d1 U6592 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][3] ), 
        .B1(n6783), .B2(\IBusCachedPlugin_cache/banks_0[1][3] ), .ZN(n6422) );
  aoi22d1 U6593 ( .A1(n6465), .A2(\IBusCachedPlugin_cache/banks_0[3][3] ), 
        .B1(n6247), .B2(\IBusCachedPlugin_cache/banks_0[7][3] ), .ZN(n6429) );
  aoi22d1 U6594 ( .A1(n6791), .A2(\IBusCachedPlugin_cache/banks_0[5][3] ), 
        .B1(n6554), .B2(\IBusCachedPlugin_cache/banks_0[4][3] ), .ZN(n6428) );
  aoi22d1 U6595 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][3] ), 
        .B1(n6696), .B2(\IBusCachedPlugin_cache/banks_0[14][3] ), .ZN(n6427)
         );
  aoi22d1 U6596 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][3] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][3] ), .ZN(n6426)
         );
  oai21d1 U6597 ( .B1(n6431), .B2(n6430), .A(n7107), .ZN(n6432) );
  oai21d1 U6598 ( .B1(n7112), .B2(n6433), .A(n6432), .ZN(n4021) );
  nd12d0 U6599 ( .A1(execute_MEMORY_ENABLE), .A2(n6996), .ZN(n4020) );
  aoi22d1 U6600 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][30] ), 
        .B1(n6784), .B2(\IBusCachedPlugin_cache/banks_0[11][30] ), .ZN(n6437)
         );
  aoi22d1 U6601 ( .A1(n6728), .A2(\IBusCachedPlugin_cache/banks_0[8][30] ), 
        .B1(n6475), .B2(\IBusCachedPlugin_cache/banks_0[12][30] ), .ZN(n6436)
         );
  aoi22d1 U6602 ( .A1(n7102), .A2(\IBusCachedPlugin_cache/banks_0[4][30] ), 
        .B1(n6696), .B2(\IBusCachedPlugin_cache/banks_0[14][30] ), .ZN(n6435)
         );
  aoi22d1 U6603 ( .A1(n6754), .A2(\IBusCachedPlugin_cache/banks_0[3][30] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][30] ), .ZN(n6434)
         );
  aoi22d1 U6604 ( .A1(n6438), .A2(\IBusCachedPlugin_cache/banks_0[10][30] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][30] ), .ZN(n6442)
         );
  aoi22d1 U6605 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][30] ), 
        .B1(n6783), .B2(\IBusCachedPlugin_cache/banks_0[1][30] ), .ZN(n6441)
         );
  aoi22d1 U6606 ( .A1(n6789), .A2(\IBusCachedPlugin_cache/banks_0[0][30] ), 
        .B1(n6637), .B2(\IBusCachedPlugin_cache/banks_0[5][30] ), .ZN(n6440)
         );
  aoi22d1 U6607 ( .A1(n6772), .A2(\IBusCachedPlugin_cache/banks_0[2][30] ), 
        .B1(n6247), .B2(\IBusCachedPlugin_cache/banks_0[7][30] ), .ZN(n6439)
         );
  oai21d1 U6608 ( .B1(n6444), .B2(n6443), .A(n7107), .ZN(n6445) );
  oai21d1 U6609 ( .B1(n7007), .B2(n6446), .A(n6445), .ZN(n4019) );
  aoi22d1 U6610 ( .A1(n6772), .A2(\IBusCachedPlugin_cache/banks_0[2][29] ), 
        .B1(n6783), .B2(\IBusCachedPlugin_cache/banks_0[1][29] ), .ZN(n6450)
         );
  aoi22d1 U6611 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][29] ), 
        .B1(n6475), .B2(\IBusCachedPlugin_cache/banks_0[12][29] ), .ZN(n6449)
         );
  aoi22d1 U6612 ( .A1(n6465), .A2(\IBusCachedPlugin_cache/banks_0[3][29] ), 
        .B1(n6784), .B2(\IBusCachedPlugin_cache/banks_0[11][29] ), .ZN(n6448)
         );
  aoi22d1 U6613 ( .A1(n6791), .A2(\IBusCachedPlugin_cache/banks_0[5][29] ), 
        .B1(n6554), .B2(\IBusCachedPlugin_cache/banks_0[4][29] ), .ZN(n6447)
         );
  aoi22d1 U6614 ( .A1(n6696), .A2(\IBusCachedPlugin_cache/banks_0[14][29] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][29] ), .ZN(n6454)
         );
  aoi22d1 U6615 ( .A1(n6789), .A2(\IBusCachedPlugin_cache/banks_0[0][29] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][29] ), .ZN(n6453)
         );
  aoi22d1 U6616 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][29] ), 
        .B1(n7097), .B2(\IBusCachedPlugin_cache/banks_0[10][29] ), .ZN(n6452)
         );
  aoi22d1 U6617 ( .A1(n6651), .A2(\IBusCachedPlugin_cache/banks_0[9][29] ), 
        .B1(n6728), .B2(\IBusCachedPlugin_cache/banks_0[8][29] ), .ZN(n6451)
         );
  oai21d1 U6618 ( .B1(n6456), .B2(n6455), .A(n7107), .ZN(n6457) );
  oai21d1 U6619 ( .B1(n7112), .B2(n6458), .A(n6457), .ZN(n4018) );
  aoim22d1 U6620 ( .A1(n6459), .A2(n7117), .B1(n6996), .B2(
        memory_INSTRUCTION_29), .Z(n4017) );
  aoi22d1 U6621 ( .A1(n6767), .A2(\IBusCachedPlugin_cache/banks_0[1][28] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][28] ), .ZN(n6464)
         );
  aoi22d1 U6622 ( .A1(n6791), .A2(\IBusCachedPlugin_cache/banks_0[5][28] ), 
        .B1(n6652), .B2(\IBusCachedPlugin_cache/banks_0[11][28] ), .ZN(n6463)
         );
  buffd1 U6623 ( .I(n6460), .Z(n7094) );
  aoi22d1 U6624 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][28] ), 
        .B1(n6554), .B2(\IBusCachedPlugin_cache/banks_0[4][28] ), .ZN(n6462)
         );
  aoi22d1 U6625 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][28] ), 
        .B1(n6772), .B2(\IBusCachedPlugin_cache/banks_0[2][28] ), .ZN(n6461)
         );
  aoi22d1 U6626 ( .A1(n6790), .A2(\IBusCachedPlugin_cache/banks_0[12][28] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][28] ), .ZN(n6469)
         );
  aoi22d1 U6627 ( .A1(n6465), .A2(\IBusCachedPlugin_cache/banks_0[3][28] ), 
        .B1(n6438), .B2(\IBusCachedPlugin_cache/banks_0[10][28] ), .ZN(n6468)
         );
  aoi22d1 U6628 ( .A1(n6537), .A2(\IBusCachedPlugin_cache/banks_0[14][28] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][28] ), .ZN(n6467)
         );
  aoi22d1 U6629 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][28] ), 
        .B1(n7095), .B2(\IBusCachedPlugin_cache/banks_0[8][28] ), .ZN(n6466)
         );
  oai21d1 U6630 ( .B1(n6471), .B2(n6470), .A(n7107), .ZN(n6472) );
  oai21d1 U6631 ( .B1(n7112), .B2(n6473), .A(n6472), .ZN(n4016) );
  aoim22d1 U6632 ( .A1(n6474), .A2(n6997), .B1(n7117), .B2(
        memory_INSTRUCTION_28), .Z(n4015) );
  aoi22d1 U6633 ( .A1(n6475), .A2(\IBusCachedPlugin_cache/banks_0[12][27] ), 
        .B1(n6696), .B2(\IBusCachedPlugin_cache/banks_0[14][27] ), .ZN(n6479)
         );
  aoi22d1 U6634 ( .A1(n6791), .A2(\IBusCachedPlugin_cache/banks_0[5][27] ), 
        .B1(n6247), .B2(\IBusCachedPlugin_cache/banks_0[7][27] ), .ZN(n6478)
         );
  aoi22d1 U6635 ( .A1(n6651), .A2(\IBusCachedPlugin_cache/banks_0[9][27] ), 
        .B1(n7102), .B2(\IBusCachedPlugin_cache/banks_0[4][27] ), .ZN(n6477)
         );
  aoi22d1 U6636 ( .A1(n6789), .A2(\IBusCachedPlugin_cache/banks_0[0][27] ), 
        .B1(n6772), .B2(\IBusCachedPlugin_cache/banks_0[2][27] ), .ZN(n6476)
         );
  aoi22d1 U6637 ( .A1(n6784), .A2(\IBusCachedPlugin_cache/banks_0[11][27] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][27] ), .ZN(n6483)
         );
  aoi22d1 U6638 ( .A1(n6754), .A2(\IBusCachedPlugin_cache/banks_0[3][27] ), 
        .B1(n6438), .B2(\IBusCachedPlugin_cache/banks_0[10][27] ), .ZN(n6482)
         );
  aoi22d1 U6639 ( .A1(n6783), .A2(\IBusCachedPlugin_cache/banks_0[1][27] ), 
        .B1(n6728), .B2(\IBusCachedPlugin_cache/banks_0[8][27] ), .ZN(n6481)
         );
  aoi22d1 U6640 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][27] ), 
        .B1(n6672), .B2(\IBusCachedPlugin_cache/banks_0[13][27] ), .ZN(n6480)
         );
  inv0d1 U6641 ( .I(n6936), .ZN(n6800) );
  oai21d1 U6642 ( .B1(n6485), .B2(n6484), .A(n6800), .ZN(n6486) );
  oai21d1 U6643 ( .B1(n7112), .B2(n6487), .A(n6486), .ZN(n4014) );
  aoi22d1 U6644 ( .A1(n7095), .A2(\IBusCachedPlugin_cache/banks_0[8][26] ), 
        .B1(n6475), .B2(\IBusCachedPlugin_cache/banks_0[12][26] ), .ZN(n6491)
         );
  aoi22d1 U6645 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][26] ), 
        .B1(n7102), .B2(\IBusCachedPlugin_cache/banks_0[4][26] ), .ZN(n6490)
         );
  aoi22d1 U6646 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][26] ), 
        .B1(n6767), .B2(\IBusCachedPlugin_cache/banks_0[1][26] ), .ZN(n6489)
         );
  aoi22d1 U6647 ( .A1(n6754), .A2(\IBusCachedPlugin_cache/banks_0[3][26] ), 
        .B1(n6247), .B2(\IBusCachedPlugin_cache/banks_0[7][26] ), .ZN(n6488)
         );
  aoi22d1 U6648 ( .A1(n7097), .A2(\IBusCachedPlugin_cache/banks_0[10][26] ), 
        .B1(n6696), .B2(\IBusCachedPlugin_cache/banks_0[14][26] ), .ZN(n6495)
         );
  aoi22d1 U6649 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][26] ), 
        .B1(n6672), .B2(\IBusCachedPlugin_cache/banks_0[13][26] ), .ZN(n6494)
         );
  aoi22d1 U6650 ( .A1(n6651), .A2(\IBusCachedPlugin_cache/banks_0[9][26] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][26] ), .ZN(n6493)
         );
  aoi22d1 U6651 ( .A1(n6637), .A2(\IBusCachedPlugin_cache/banks_0[5][26] ), 
        .B1(n6652), .B2(\IBusCachedPlugin_cache/banks_0[11][26] ), .ZN(n6492)
         );
  oai21d1 U6652 ( .B1(n6497), .B2(n6496), .A(n6800), .ZN(n6498) );
  oai21d1 U6653 ( .B1(n7112), .B2(n6499), .A(n6498), .ZN(n4013) );
  aoi22d1 U6654 ( .A1(n6767), .A2(\IBusCachedPlugin_cache/banks_0[1][25] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][25] ), .ZN(n6503)
         );
  aoi22d1 U6655 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][25] ), 
        .B1(n6672), .B2(\IBusCachedPlugin_cache/banks_0[13][25] ), .ZN(n6502)
         );
  aoi22d1 U6656 ( .A1(n6772), .A2(\IBusCachedPlugin_cache/banks_0[2][25] ), 
        .B1(n6728), .B2(\IBusCachedPlugin_cache/banks_0[8][25] ), .ZN(n6501)
         );
  aoi22d1 U6657 ( .A1(n6784), .A2(\IBusCachedPlugin_cache/banks_0[11][25] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][25] ), .ZN(n6500)
         );
  aoi22d1 U6658 ( .A1(n6791), .A2(\IBusCachedPlugin_cache/banks_0[5][25] ), 
        .B1(n7102), .B2(\IBusCachedPlugin_cache/banks_0[4][25] ), .ZN(n6507)
         );
  aoi22d1 U6659 ( .A1(n6754), .A2(\IBusCachedPlugin_cache/banks_0[3][25] ), 
        .B1(n7097), .B2(\IBusCachedPlugin_cache/banks_0[10][25] ), .ZN(n6506)
         );
  aoi22d1 U6660 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][25] ), 
        .B1(n6696), .B2(\IBusCachedPlugin_cache/banks_0[14][25] ), .ZN(n6505)
         );
  aoi22d1 U6661 ( .A1(n6790), .A2(\IBusCachedPlugin_cache/banks_0[12][25] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][25] ), .ZN(n6504)
         );
  oai21d1 U6662 ( .B1(n6509), .B2(n6508), .A(n6800), .ZN(n6510) );
  oai21d1 U6663 ( .B1(n7112), .B2(n6511), .A(n6510), .ZN(n4012) );
  aoi22d1 U6664 ( .A1(n6754), .A2(\IBusCachedPlugin_cache/banks_0[3][24] ), 
        .B1(n6767), .B2(\IBusCachedPlugin_cache/banks_0[1][24] ), .ZN(n6515)
         );
  aoi22d1 U6665 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][24] ), 
        .B1(n6772), .B2(\IBusCachedPlugin_cache/banks_0[2][24] ), .ZN(n6514)
         );
  aoi22d1 U6666 ( .A1(n6652), .A2(\IBusCachedPlugin_cache/banks_0[11][24] ), 
        .B1(n6696), .B2(\IBusCachedPlugin_cache/banks_0[14][24] ), .ZN(n6513)
         );
  aoi22d1 U6667 ( .A1(n7097), .A2(\IBusCachedPlugin_cache/banks_0[10][24] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][24] ), .ZN(n6512)
         );
  aoi22d1 U6668 ( .A1(n6789), .A2(\IBusCachedPlugin_cache/banks_0[0][24] ), 
        .B1(n6637), .B2(\IBusCachedPlugin_cache/banks_0[5][24] ), .ZN(n6519)
         );
  aoi22d1 U6669 ( .A1(n6651), .A2(\IBusCachedPlugin_cache/banks_0[9][24] ), 
        .B1(n6671), .B2(\IBusCachedPlugin_cache/banks_0[15][24] ), .ZN(n6518)
         );
  aoi22d1 U6670 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][24] ), 
        .B1(n6475), .B2(\IBusCachedPlugin_cache/banks_0[12][24] ), .ZN(n6517)
         );
  aoi22d1 U6671 ( .A1(n6554), .A2(\IBusCachedPlugin_cache/banks_0[4][24] ), 
        .B1(n6728), .B2(\IBusCachedPlugin_cache/banks_0[8][24] ), .ZN(n6516)
         );
  oai21d1 U6672 ( .B1(n6521), .B2(n6520), .A(n6800), .ZN(n6522) );
  oai21d1 U6673 ( .B1(n7112), .B2(n6523), .A(n6522), .ZN(n4011) );
  aoi22d1 U6674 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][23] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][23] ), .ZN(n6527)
         );
  aoi22d1 U6675 ( .A1(n6637), .A2(\IBusCachedPlugin_cache/banks_0[5][23] ), 
        .B1(n7102), .B2(\IBusCachedPlugin_cache/banks_0[4][23] ), .ZN(n6526)
         );
  aoi22d1 U6676 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][23] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][23] ), .ZN(n6525)
         );
  aoi22d1 U6677 ( .A1(n7097), .A2(\IBusCachedPlugin_cache/banks_0[10][23] ), 
        .B1(n6696), .B2(\IBusCachedPlugin_cache/banks_0[14][23] ), .ZN(n6524)
         );
  aoi22d1 U6678 ( .A1(n6528), .A2(\IBusCachedPlugin_cache/banks_0[8][23] ), 
        .B1(n6475), .B2(\IBusCachedPlugin_cache/banks_0[12][23] ), .ZN(n6532)
         );
  aoi22d1 U6679 ( .A1(n6767), .A2(\IBusCachedPlugin_cache/banks_0[1][23] ), 
        .B1(n6652), .B2(\IBusCachedPlugin_cache/banks_0[11][23] ), .ZN(n6531)
         );
  aoi22d1 U6680 ( .A1(n6789), .A2(\IBusCachedPlugin_cache/banks_0[0][23] ), 
        .B1(n6772), .B2(\IBusCachedPlugin_cache/banks_0[2][23] ), .ZN(n6530)
         );
  aoi22d1 U6681 ( .A1(n6465), .A2(\IBusCachedPlugin_cache/banks_0[3][23] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][23] ), .ZN(n6529)
         );
  oai21d1 U6682 ( .B1(n6534), .B2(n6533), .A(n6800), .ZN(n6535) );
  oai21d1 U6683 ( .B1(n7112), .B2(n6536), .A(n6535), .ZN(n4010) );
  aoi22d1 U6684 ( .A1(n6772), .A2(\IBusCachedPlugin_cache/banks_0[2][22] ), 
        .B1(n7097), .B2(\IBusCachedPlugin_cache/banks_0[10][22] ), .ZN(n6541)
         );
  aoi22d1 U6685 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][22] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][22] ), .ZN(n6540)
         );
  aoi22d1 U6686 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][22] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][22] ), .ZN(n6539)
         );
  aoi22d1 U6687 ( .A1(n6537), .A2(\IBusCachedPlugin_cache/banks_0[14][22] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][22] ), .ZN(n6538)
         );
  aoi22d1 U6688 ( .A1(n6465), .A2(\IBusCachedPlugin_cache/banks_0[3][22] ), 
        .B1(n6790), .B2(\IBusCachedPlugin_cache/banks_0[12][22] ), .ZN(n6545)
         );
  aoi22d1 U6689 ( .A1(n6783), .A2(\IBusCachedPlugin_cache/banks_0[1][22] ), 
        .B1(n6728), .B2(\IBusCachedPlugin_cache/banks_0[8][22] ), .ZN(n6544)
         );
  aoi22d1 U6690 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][22] ), 
        .B1(n6652), .B2(\IBusCachedPlugin_cache/banks_0[11][22] ), .ZN(n6543)
         );
  aoi22d1 U6691 ( .A1(n6637), .A2(\IBusCachedPlugin_cache/banks_0[5][22] ), 
        .B1(n7102), .B2(\IBusCachedPlugin_cache/banks_0[4][22] ), .ZN(n6542)
         );
  oai21d1 U6692 ( .B1(n6547), .B2(n6546), .A(n6800), .ZN(n6548) );
  oai21d1 U6693 ( .B1(n7112), .B2(n6549), .A(n6548), .ZN(n4009) );
  aoi22d1 U6694 ( .A1(n6772), .A2(\IBusCachedPlugin_cache/banks_0[2][21] ), 
        .B1(n6696), .B2(\IBusCachedPlugin_cache/banks_0[14][21] ), .ZN(n6553)
         );
  aoi22d1 U6695 ( .A1(n6465), .A2(\IBusCachedPlugin_cache/banks_0[3][21] ), 
        .B1(n6784), .B2(\IBusCachedPlugin_cache/banks_0[11][21] ), .ZN(n6552)
         );
  aoi22d1 U6696 ( .A1(n6767), .A2(\IBusCachedPlugin_cache/banks_0[1][21] ), 
        .B1(n6728), .B2(\IBusCachedPlugin_cache/banks_0[8][21] ), .ZN(n6551)
         );
  aoi22d1 U6697 ( .A1(n6791), .A2(\IBusCachedPlugin_cache/banks_0[5][21] ), 
        .B1(n6672), .B2(\IBusCachedPlugin_cache/banks_0[13][21] ), .ZN(n6550)
         );
  aoi22d1 U6698 ( .A1(n7097), .A2(\IBusCachedPlugin_cache/banks_0[10][21] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][21] ), .ZN(n6558)
         );
  aoi22d1 U6699 ( .A1(n6651), .A2(\IBusCachedPlugin_cache/banks_0[9][21] ), 
        .B1(n6790), .B2(\IBusCachedPlugin_cache/banks_0[12][21] ), .ZN(n6557)
         );
  aoi22d1 U6700 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][21] ), 
        .B1(n6789), .B2(\IBusCachedPlugin_cache/banks_0[0][21] ), .ZN(n6556)
         );
  aoi22d1 U6701 ( .A1(n6554), .A2(\IBusCachedPlugin_cache/banks_0[4][21] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][21] ), .ZN(n6555)
         );
  oai21d1 U6702 ( .B1(n6560), .B2(n6559), .A(n6800), .ZN(n6561) );
  oai21d1 U6703 ( .B1(n7112), .B2(n6562), .A(n6561), .ZN(n4008) );
  aoi22d1 U6704 ( .A1(n6628), .A2(\IBusCachedPlugin_cache/banks_0[6][20] ), 
        .B1(n6438), .B2(\IBusCachedPlugin_cache/banks_0[10][20] ), .ZN(n6566)
         );
  aoi22d1 U6705 ( .A1(n6652), .A2(\IBusCachedPlugin_cache/banks_0[11][20] ), 
        .B1(n6728), .B2(\IBusCachedPlugin_cache/banks_0[8][20] ), .ZN(n6565)
         );
  aoi22d1 U6706 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][20] ), 
        .B1(n6791), .B2(\IBusCachedPlugin_cache/banks_0[5][20] ), .ZN(n6564)
         );
  aoi22d1 U6707 ( .A1(n6465), .A2(\IBusCachedPlugin_cache/banks_0[3][20] ), 
        .B1(n6767), .B2(\IBusCachedPlugin_cache/banks_0[1][20] ), .ZN(n6563)
         );
  aoi22d1 U6708 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][20] ), 
        .B1(n6672), .B2(\IBusCachedPlugin_cache/banks_0[13][20] ), .ZN(n6570)
         );
  aoi22d1 U6709 ( .A1(n6537), .A2(\IBusCachedPlugin_cache/banks_0[14][20] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][20] ), .ZN(n6569)
         );
  aoi22d1 U6710 ( .A1(n6790), .A2(\IBusCachedPlugin_cache/banks_0[12][20] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][20] ), .ZN(n6568)
         );
  aoi22d1 U6711 ( .A1(n6651), .A2(\IBusCachedPlugin_cache/banks_0[9][20] ), 
        .B1(n7102), .B2(\IBusCachedPlugin_cache/banks_0[4][20] ), .ZN(n6567)
         );
  oai21d1 U6712 ( .B1(n6572), .B2(n6571), .A(n6800), .ZN(n6573) );
  oai21d1 U6713 ( .B1(n7112), .B2(n6574), .A(n6573), .ZN(n4007) );
  aoi22d1 U6714 ( .A1(n6554), .A2(\IBusCachedPlugin_cache/banks_0[4][19] ), 
        .B1(n6475), .B2(\IBusCachedPlugin_cache/banks_0[12][19] ), .ZN(n6578)
         );
  aoi22d1 U6715 ( .A1(n7095), .A2(\IBusCachedPlugin_cache/banks_0[8][19] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][19] ), .ZN(n6577)
         );
  aoi22d1 U6716 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][19] ), 
        .B1(n6754), .B2(\IBusCachedPlugin_cache/banks_0[3][19] ), .ZN(n6576)
         );
  aoi22d1 U6717 ( .A1(n6651), .A2(\IBusCachedPlugin_cache/banks_0[9][19] ), 
        .B1(n6696), .B2(\IBusCachedPlugin_cache/banks_0[14][19] ), .ZN(n6575)
         );
  aoi22d1 U6718 ( .A1(n7097), .A2(\IBusCachedPlugin_cache/banks_0[10][19] ), 
        .B1(n6671), .B2(\IBusCachedPlugin_cache/banks_0[15][19] ), .ZN(n6582)
         );
  aoi22d1 U6719 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][19] ), 
        .B1(n6652), .B2(\IBusCachedPlugin_cache/banks_0[11][19] ), .ZN(n6581)
         );
  aoi22d1 U6720 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][19] ), 
        .B1(n6767), .B2(\IBusCachedPlugin_cache/banks_0[1][19] ), .ZN(n6580)
         );
  aoi22d1 U6721 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][19] ), 
        .B1(n6637), .B2(\IBusCachedPlugin_cache/banks_0[5][19] ), .ZN(n6579)
         );
  oai21d1 U6722 ( .B1(n6584), .B2(n6583), .A(n6800), .ZN(n6585) );
  oai21d1 U6723 ( .B1(n7112), .B2(n6586), .A(n6585), .ZN(n4006) );
  aoi22d1 U6724 ( .A1(n6783), .A2(\IBusCachedPlugin_cache/banks_0[1][18] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][18] ), .ZN(n6590)
         );
  aoi22d1 U6725 ( .A1(n7102), .A2(\IBusCachedPlugin_cache/banks_0[4][18] ), 
        .B1(n6728), .B2(\IBusCachedPlugin_cache/banks_0[8][18] ), .ZN(n6589)
         );
  aoi22d1 U6726 ( .A1(n6537), .A2(\IBusCachedPlugin_cache/banks_0[14][18] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][18] ), .ZN(n6588)
         );
  aoi22d1 U6727 ( .A1(n6637), .A2(\IBusCachedPlugin_cache/banks_0[5][18] ), 
        .B1(n6672), .B2(\IBusCachedPlugin_cache/banks_0[13][18] ), .ZN(n6587)
         );
  aoi22d1 U6728 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][18] ), 
        .B1(n6789), .B2(\IBusCachedPlugin_cache/banks_0[0][18] ), .ZN(n6594)
         );
  aoi22d1 U6729 ( .A1(n6465), .A2(\IBusCachedPlugin_cache/banks_0[3][18] ), 
        .B1(n6652), .B2(\IBusCachedPlugin_cache/banks_0[11][18] ), .ZN(n6593)
         );
  aoi22d1 U6730 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][18] ), 
        .B1(n6438), .B2(\IBusCachedPlugin_cache/banks_0[10][18] ), .ZN(n6592)
         );
  aoi22d1 U6731 ( .A1(n6790), .A2(\IBusCachedPlugin_cache/banks_0[12][18] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][18] ), .ZN(n6591)
         );
  oai21d1 U6732 ( .B1(n6596), .B2(n6595), .A(n2356), .ZN(n6597) );
  oai21d1 U6733 ( .B1(n7112), .B2(n6598), .A(n6597), .ZN(n4005) );
  aoi22d1 U6734 ( .A1(n6599), .A2(\IBusCachedPlugin_cache/banks_0[6][17] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][17] ), .ZN(n6603)
         );
  aoi22d1 U6735 ( .A1(n6790), .A2(\IBusCachedPlugin_cache/banks_0[12][17] ), 
        .B1(n6671), .B2(\IBusCachedPlugin_cache/banks_0[15][17] ), .ZN(n6602)
         );
  aoi22d1 U6736 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][17] ), 
        .B1(n6791), .B2(\IBusCachedPlugin_cache/banks_0[5][17] ), .ZN(n6601)
         );
  aoi22d1 U6737 ( .A1(n6465), .A2(\IBusCachedPlugin_cache/banks_0[3][17] ), 
        .B1(n6728), .B2(\IBusCachedPlugin_cache/banks_0[8][17] ), .ZN(n6600)
         );
  aoi22d1 U6738 ( .A1(n6783), .A2(\IBusCachedPlugin_cache/banks_0[1][17] ), 
        .B1(n6696), .B2(\IBusCachedPlugin_cache/banks_0[14][17] ), .ZN(n6607)
         );
  aoi22d1 U6739 ( .A1(n6438), .A2(\IBusCachedPlugin_cache/banks_0[10][17] ), 
        .B1(n7102), .B2(\IBusCachedPlugin_cache/banks_0[4][17] ), .ZN(n6606)
         );
  aoi22d1 U6740 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][17] ), 
        .B1(n6652), .B2(\IBusCachedPlugin_cache/banks_0[11][17] ), .ZN(n6605)
         );
  aoi22d1 U6741 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][17] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][17] ), .ZN(n6604)
         );
  oai21d1 U6742 ( .B1(n6609), .B2(n6608), .A(n6800), .ZN(n6610) );
  oai21d1 U6743 ( .B1(n7112), .B2(n6611), .A(n6610), .ZN(n4004) );
  aoi22d1 U6744 ( .A1(n6784), .A2(\IBusCachedPlugin_cache/banks_0[11][16] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][16] ), .ZN(n6615)
         );
  aoi22d1 U6745 ( .A1(n6767), .A2(\IBusCachedPlugin_cache/banks_0[1][16] ), 
        .B1(n7102), .B2(\IBusCachedPlugin_cache/banks_0[4][16] ), .ZN(n6614)
         );
  aoi22d1 U6746 ( .A1(n6628), .A2(\IBusCachedPlugin_cache/banks_0[6][16] ), 
        .B1(n6672), .B2(\IBusCachedPlugin_cache/banks_0[13][16] ), .ZN(n6613)
         );
  aoi22d1 U6747 ( .A1(n6637), .A2(\IBusCachedPlugin_cache/banks_0[5][16] ), 
        .B1(n6475), .B2(\IBusCachedPlugin_cache/banks_0[12][16] ), .ZN(n6612)
         );
  aoi22d1 U6748 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][16] ), 
        .B1(n7095), .B2(\IBusCachedPlugin_cache/banks_0[8][16] ), .ZN(n6619)
         );
  aoi22d1 U6749 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][16] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][16] ), .ZN(n6618)
         );
  aoi22d1 U6750 ( .A1(n6465), .A2(\IBusCachedPlugin_cache/banks_0[3][16] ), 
        .B1(n7097), .B2(\IBusCachedPlugin_cache/banks_0[10][16] ), .ZN(n6617)
         );
  aoi22d1 U6751 ( .A1(n6696), .A2(\IBusCachedPlugin_cache/banks_0[14][16] ), 
        .B1(n6671), .B2(\IBusCachedPlugin_cache/banks_0[15][16] ), .ZN(n6616)
         );
  oai21d1 U6752 ( .B1(n6621), .B2(n6620), .A(n2356), .ZN(n6622) );
  oai21d1 U6753 ( .B1(n7112), .B2(n6623), .A(n6622), .ZN(n4003) );
  aoi22d1 U6754 ( .A1(n6537), .A2(\IBusCachedPlugin_cache/banks_0[14][15] ), 
        .B1(n6247), .B2(\IBusCachedPlugin_cache/banks_0[7][15] ), .ZN(n6627)
         );
  aoi22d1 U6755 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][15] ), 
        .B1(n6728), .B2(\IBusCachedPlugin_cache/banks_0[8][15] ), .ZN(n6626)
         );
  aoi22d1 U6756 ( .A1(n6465), .A2(\IBusCachedPlugin_cache/banks_0[3][15] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][15] ), .ZN(n6625)
         );
  aoi22d1 U6757 ( .A1(n6637), .A2(\IBusCachedPlugin_cache/banks_0[5][15] ), 
        .B1(n6475), .B2(\IBusCachedPlugin_cache/banks_0[12][15] ), .ZN(n6624)
         );
  aoi22d1 U6758 ( .A1(n6628), .A2(\IBusCachedPlugin_cache/banks_0[6][15] ), 
        .B1(n7102), .B2(\IBusCachedPlugin_cache/banks_0[4][15] ), .ZN(n6632)
         );
  aoi22d1 U6759 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][15] ), 
        .B1(n6671), .B2(\IBusCachedPlugin_cache/banks_0[15][15] ), .ZN(n6631)
         );
  aoi22d1 U6760 ( .A1(n6438), .A2(\IBusCachedPlugin_cache/banks_0[10][15] ), 
        .B1(n6784), .B2(\IBusCachedPlugin_cache/banks_0[11][15] ), .ZN(n6630)
         );
  aoi22d1 U6761 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][15] ), 
        .B1(n6767), .B2(\IBusCachedPlugin_cache/banks_0[1][15] ), .ZN(n6629)
         );
  oai21d1 U6762 ( .B1(n6634), .B2(n6633), .A(n2356), .ZN(n6635) );
  oai21d1 U6763 ( .B1(n7112), .B2(n6636), .A(n6635), .ZN(n4002) );
  aoi22d1 U6764 ( .A1(n6790), .A2(\IBusCachedPlugin_cache/banks_0[12][14] ), 
        .B1(n6247), .B2(\IBusCachedPlugin_cache/banks_0[7][14] ), .ZN(n6641)
         );
  aoi22d1 U6765 ( .A1(n6637), .A2(\IBusCachedPlugin_cache/banks_0[5][14] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][14] ), .ZN(n6640)
         );
  aoi22d1 U6766 ( .A1(n7102), .A2(\IBusCachedPlugin_cache/banks_0[4][14] ), 
        .B1(n6696), .B2(\IBusCachedPlugin_cache/banks_0[14][14] ), .ZN(n6639)
         );
  aoi22d1 U6767 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][14] ), 
        .B1(n6767), .B2(\IBusCachedPlugin_cache/banks_0[1][14] ), .ZN(n6638)
         );
  aoi22d1 U6768 ( .A1(n6628), .A2(\IBusCachedPlugin_cache/banks_0[6][14] ), 
        .B1(n7095), .B2(\IBusCachedPlugin_cache/banks_0[8][14] ), .ZN(n6645)
         );
  aoi22d1 U6769 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][14] ), 
        .B1(n6438), .B2(\IBusCachedPlugin_cache/banks_0[10][14] ), .ZN(n6644)
         );
  aoi22d1 U6770 ( .A1(n6784), .A2(\IBusCachedPlugin_cache/banks_0[11][14] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][14] ), .ZN(n6643)
         );
  aoi22d1 U6771 ( .A1(n6465), .A2(\IBusCachedPlugin_cache/banks_0[3][14] ), 
        .B1(n6672), .B2(\IBusCachedPlugin_cache/banks_0[13][14] ), .ZN(n6642)
         );
  oai21d1 U6772 ( .B1(n6647), .B2(n6646), .A(n7085), .ZN(n6648) );
  oai21d1 U6773 ( .B1(n7112), .B2(n6649), .A(n6648), .ZN(n4001) );
  aoim22d1 U6774 ( .A1(n6650), .A2(n6996), .B1(n6996), .B2(
        memory_INSTRUCTION[14]), .Z(n4000) );
  aoi22d1 U6775 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][13] ), 
        .B1(n6791), .B2(\IBusCachedPlugin_cache/banks_0[5][13] ), .ZN(n6656)
         );
  aoi22d1 U6776 ( .A1(n6651), .A2(\IBusCachedPlugin_cache/banks_0[9][13] ), 
        .B1(n7102), .B2(\IBusCachedPlugin_cache/banks_0[4][13] ), .ZN(n6655)
         );
  aoi22d1 U6777 ( .A1(n6652), .A2(\IBusCachedPlugin_cache/banks_0[11][13] ), 
        .B1(n6671), .B2(\IBusCachedPlugin_cache/banks_0[15][13] ), .ZN(n6654)
         );
  aoi22d1 U6778 ( .A1(n6628), .A2(\IBusCachedPlugin_cache/banks_0[6][13] ), 
        .B1(n6475), .B2(\IBusCachedPlugin_cache/banks_0[12][13] ), .ZN(n6653)
         );
  aoi22d1 U6779 ( .A1(n6438), .A2(\IBusCachedPlugin_cache/banks_0[10][13] ), 
        .B1(n6537), .B2(\IBusCachedPlugin_cache/banks_0[14][13] ), .ZN(n6660)
         );
  aoi22d1 U6780 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][13] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][13] ), .ZN(n6659)
         );
  aoi22d1 U6781 ( .A1(n6754), .A2(\IBusCachedPlugin_cache/banks_0[3][13] ), 
        .B1(n6767), .B2(\IBusCachedPlugin_cache/banks_0[1][13] ), .ZN(n6658)
         );
  aoi22d1 U6782 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][13] ), 
        .B1(n6728), .B2(\IBusCachedPlugin_cache/banks_0[8][13] ), .ZN(n6657)
         );
  oai21d1 U6783 ( .B1(n6662), .B2(n6661), .A(n2356), .ZN(n6663) );
  oai21d1 U6784 ( .B1(n6800), .B2(n6664), .A(n6663), .ZN(n3999) );
  nr02d1 U6785 ( .A1(n6977), .A2(n6919), .ZN(n6988) );
  inv0d0 U6786 ( .I(n6988), .ZN(n6986) );
  oai21d1 U6787 ( .B1(n6993), .B2(n6665), .A(n6986), .ZN(n3998) );
  aoim22d1 U6788 ( .A1(n6666), .A2(n6997), .B1(n6997), .B2(
        memory_INSTRUCTION[13]), .Z(n3997) );
  aoi22d1 U6789 ( .A1(n6791), .A2(\IBusCachedPlugin_cache/banks_0[5][12] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][12] ), .ZN(n6670)
         );
  aoi22d1 U6790 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][12] ), 
        .B1(n6754), .B2(\IBusCachedPlugin_cache/banks_0[3][12] ), .ZN(n6669)
         );
  aoi22d1 U6791 ( .A1(n6628), .A2(\IBusCachedPlugin_cache/banks_0[6][12] ), 
        .B1(n6554), .B2(\IBusCachedPlugin_cache/banks_0[4][12] ), .ZN(n6668)
         );
  aoi22d1 U6792 ( .A1(n7095), .A2(\IBusCachedPlugin_cache/banks_0[8][12] ), 
        .B1(n6537), .B2(\IBusCachedPlugin_cache/banks_0[14][12] ), .ZN(n6667)
         );
  aoi22d1 U6793 ( .A1(n6438), .A2(\IBusCachedPlugin_cache/banks_0[10][12] ), 
        .B1(n6783), .B2(\IBusCachedPlugin_cache/banks_0[1][12] ), .ZN(n6676)
         );
  aoi22d1 U6794 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][12] ), 
        .B1(n6671), .B2(\IBusCachedPlugin_cache/banks_0[15][12] ), .ZN(n6675)
         );
  aoi22d1 U6795 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][12] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][12] ), .ZN(n6674)
         );
  aoi22d1 U6796 ( .A1(n6652), .A2(\IBusCachedPlugin_cache/banks_0[11][12] ), 
        .B1(n6790), .B2(\IBusCachedPlugin_cache/banks_0[12][12] ), .ZN(n6673)
         );
  oai21d1 U6797 ( .B1(n6678), .B2(n6677), .A(n2356), .ZN(n6679) );
  oai21d1 U6798 ( .B1(n7107), .B2(n6680), .A(n6679), .ZN(n3996) );
  aoim22d1 U6799 ( .A1(n6681), .A2(n6996), .B1(n6996), .B2(
        memory_INSTRUCTION[12]), .Z(n3995) );
  aoim22d1 U6800 ( .A1(n6681), .A2(n6972), .B1(n6993), .B2(
        dBus_cmd_halfPipe_payload_size[0]), .Z(n3994) );
  aoi22d1 U6801 ( .A1(n6754), .A2(\IBusCachedPlugin_cache/banks_0[3][11] ), 
        .B1(n6672), .B2(\IBusCachedPlugin_cache/banks_0[13][11] ), .ZN(n6685)
         );
  aoi22d1 U6802 ( .A1(n6790), .A2(\IBusCachedPlugin_cache/banks_0[12][11] ), 
        .B1(n6671), .B2(\IBusCachedPlugin_cache/banks_0[15][11] ), .ZN(n6684)
         );
  aoi22d1 U6803 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][11] ), 
        .B1(n6554), .B2(\IBusCachedPlugin_cache/banks_0[4][11] ), .ZN(n6683)
         );
  aoi22d1 U6804 ( .A1(n6789), .A2(\IBusCachedPlugin_cache/banks_0[0][11] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][11] ), .ZN(n6682)
         );
  aoi22d1 U6805 ( .A1(n6537), .A2(\IBusCachedPlugin_cache/banks_0[14][11] ), 
        .B1(n6247), .B2(\IBusCachedPlugin_cache/banks_0[7][11] ), .ZN(n6689)
         );
  aoi22d1 U6806 ( .A1(n6628), .A2(\IBusCachedPlugin_cache/banks_0[6][11] ), 
        .B1(n6783), .B2(\IBusCachedPlugin_cache/banks_0[1][11] ), .ZN(n6688)
         );
  aoi22d1 U6807 ( .A1(n6791), .A2(\IBusCachedPlugin_cache/banks_0[5][11] ), 
        .B1(n6652), .B2(\IBusCachedPlugin_cache/banks_0[11][11] ), .ZN(n6687)
         );
  aoi22d1 U6808 ( .A1(n7097), .A2(\IBusCachedPlugin_cache/banks_0[10][11] ), 
        .B1(n7095), .B2(\IBusCachedPlugin_cache/banks_0[8][11] ), .ZN(n6686)
         );
  oai21d1 U6809 ( .B1(n6691), .B2(n6690), .A(n2356), .ZN(n6692) );
  oai21d1 U6810 ( .B1(n7107), .B2(n6693), .A(n6692), .ZN(n3993) );
  aoi22d1 U6811 ( .A1(n6740), .A2(n6695), .B1(n6694), .B2(n6997), .ZN(n3992)
         );
  aoi22d1 U6812 ( .A1(n6772), .A2(\IBusCachedPlugin_cache/banks_0[2][10] ), 
        .B1(n6696), .B2(\IBusCachedPlugin_cache/banks_0[14][10] ), .ZN(n6700)
         );
  aoi22d1 U6813 ( .A1(n6791), .A2(\IBusCachedPlugin_cache/banks_0[5][10] ), 
        .B1(n6672), .B2(\IBusCachedPlugin_cache/banks_0[13][10] ), .ZN(n6699)
         );
  aoi22d1 U6814 ( .A1(n6754), .A2(\IBusCachedPlugin_cache/banks_0[3][10] ), 
        .B1(n6767), .B2(\IBusCachedPlugin_cache/banks_0[1][10] ), .ZN(n6698)
         );
  aoi22d1 U6815 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][10] ), 
        .B1(n6247), .B2(\IBusCachedPlugin_cache/banks_0[7][10] ), .ZN(n6697)
         );
  aoi22d1 U6816 ( .A1(n7102), .A2(\IBusCachedPlugin_cache/banks_0[4][10] ), 
        .B1(n6671), .B2(\IBusCachedPlugin_cache/banks_0[15][10] ), .ZN(n6704)
         );
  aoi22d1 U6817 ( .A1(n6438), .A2(\IBusCachedPlugin_cache/banks_0[10][10] ), 
        .B1(n6784), .B2(\IBusCachedPlugin_cache/banks_0[11][10] ), .ZN(n6703)
         );
  aoi22d1 U6818 ( .A1(n6628), .A2(\IBusCachedPlugin_cache/banks_0[6][10] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][10] ), .ZN(n6702)
         );
  aoi22d1 U6819 ( .A1(n6728), .A2(\IBusCachedPlugin_cache/banks_0[8][10] ), 
        .B1(n6790), .B2(\IBusCachedPlugin_cache/banks_0[12][10] ), .ZN(n6701)
         );
  oai21d1 U6820 ( .B1(n6706), .B2(n6705), .A(n2356), .ZN(n6707) );
  oai21d1 U6821 ( .B1(n7107), .B2(n6708), .A(n6707), .ZN(n3991) );
  aoim22d1 U6822 ( .A1(n6709), .A2(n6997), .B1(n7117), .B2(
        memory_INSTRUCTION[10]), .Z(n3990) );
  aoi22d1 U6823 ( .A1(n6728), .A2(\IBusCachedPlugin_cache/banks_0[8][9] ), 
        .B1(n6475), .B2(\IBusCachedPlugin_cache/banks_0[12][9] ), .ZN(n6713)
         );
  aoi22d1 U6824 ( .A1(n6628), .A2(\IBusCachedPlugin_cache/banks_0[6][9] ), 
        .B1(n6783), .B2(\IBusCachedPlugin_cache/banks_0[1][9] ), .ZN(n6712) );
  aoi22d1 U6825 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][9] ), 
        .B1(n6754), .B2(\IBusCachedPlugin_cache/banks_0[3][9] ), .ZN(n6711) );
  aoi22d1 U6826 ( .A1(n6784), .A2(\IBusCachedPlugin_cache/banks_0[11][9] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][9] ), .ZN(n6710) );
  aoi22d1 U6827 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][9] ), 
        .B1(n6637), .B2(\IBusCachedPlugin_cache/banks_0[5][9] ), .ZN(n6717) );
  aoi22d1 U6828 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][9] ), 
        .B1(n6438), .B2(\IBusCachedPlugin_cache/banks_0[10][9] ), .ZN(n6716)
         );
  aoi22d1 U6829 ( .A1(n6554), .A2(\IBusCachedPlugin_cache/banks_0[4][9] ), 
        .B1(n6671), .B2(\IBusCachedPlugin_cache/banks_0[15][9] ), .ZN(n6715)
         );
  aoi22d1 U6830 ( .A1(n6651), .A2(\IBusCachedPlugin_cache/banks_0[9][9] ), 
        .B1(n6537), .B2(\IBusCachedPlugin_cache/banks_0[14][9] ), .ZN(n6714)
         );
  oai21d1 U6831 ( .B1(n6719), .B2(n6718), .A(n2356), .ZN(n6720) );
  oai21d1 U6832 ( .B1(n6800), .B2(n6721), .A(n6720), .ZN(n3989) );
  aoim22d1 U6833 ( .A1(n6722), .A2(n6997), .B1(n6997), .B2(
        memory_INSTRUCTION[9]), .Z(n3988) );
  aoi22d1 U6834 ( .A1(n6754), .A2(\IBusCachedPlugin_cache/banks_0[3][8] ), 
        .B1(n6790), .B2(\IBusCachedPlugin_cache/banks_0[12][8] ), .ZN(n6727)
         );
  aoi22d1 U6835 ( .A1(n6637), .A2(\IBusCachedPlugin_cache/banks_0[5][8] ), 
        .B1(n6723), .B2(\IBusCachedPlugin_cache/banks_0[7][8] ), .ZN(n6726) );
  aoi22d1 U6836 ( .A1(n6652), .A2(\IBusCachedPlugin_cache/banks_0[11][8] ), 
        .B1(n6537), .B2(\IBusCachedPlugin_cache/banks_0[14][8] ), .ZN(n6725)
         );
  aoi22d1 U6837 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][8] ), 
        .B1(n6438), .B2(\IBusCachedPlugin_cache/banks_0[10][8] ), .ZN(n6724)
         );
  aoi22d1 U6838 ( .A1(n6651), .A2(\IBusCachedPlugin_cache/banks_0[9][8] ), 
        .B1(n6554), .B2(\IBusCachedPlugin_cache/banks_0[4][8] ), .ZN(n6733) );
  aoi22d1 U6839 ( .A1(n6628), .A2(\IBusCachedPlugin_cache/banks_0[6][8] ), 
        .B1(n6728), .B2(\IBusCachedPlugin_cache/banks_0[8][8] ), .ZN(n6732) );
  aoi22d1 U6840 ( .A1(n6783), .A2(\IBusCachedPlugin_cache/banks_0[1][8] ), 
        .B1(n6729), .B2(\IBusCachedPlugin_cache/banks_0[15][8] ), .ZN(n6731)
         );
  aoi22d1 U6841 ( .A1(n6789), .A2(\IBusCachedPlugin_cache/banks_0[0][8] ), 
        .B1(n6772), .B2(\IBusCachedPlugin_cache/banks_0[2][8] ), .ZN(n6730) );
  oai21d1 U6842 ( .B1(n6735), .B2(n6734), .A(n2356), .ZN(n6736) );
  oai21d1 U6843 ( .B1(n7107), .B2(n6737), .A(n6736), .ZN(n3987) );
  aoi22d1 U6844 ( .A1(n6740), .A2(n6739), .B1(n6738), .B2(n7117), .ZN(n3986)
         );
  aoi22d1 U6845 ( .A1(n6475), .A2(\IBusCachedPlugin_cache/banks_0[12][7] ), 
        .B1(n6671), .B2(\IBusCachedPlugin_cache/banks_0[15][7] ), .ZN(n6744)
         );
  aoi22d1 U6846 ( .A1(n6628), .A2(\IBusCachedPlugin_cache/banks_0[6][7] ), 
        .B1(n7095), .B2(\IBusCachedPlugin_cache/banks_0[8][7] ), .ZN(n6743) );
  aoi22d1 U6847 ( .A1(n6438), .A2(\IBusCachedPlugin_cache/banks_0[10][7] ), 
        .B1(n6554), .B2(\IBusCachedPlugin_cache/banks_0[4][7] ), .ZN(n6742) );
  aoi22d1 U6848 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][7] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][7] ), .ZN(n6741) );
  aoi22d1 U6849 ( .A1(n6789), .A2(\IBusCachedPlugin_cache/banks_0[0][7] ), 
        .B1(n6783), .B2(\IBusCachedPlugin_cache/banks_0[1][7] ), .ZN(n6748) );
  aoi22d1 U6850 ( .A1(n6537), .A2(\IBusCachedPlugin_cache/banks_0[14][7] ), 
        .B1(n6247), .B2(\IBusCachedPlugin_cache/banks_0[7][7] ), .ZN(n6747) );
  aoi22d1 U6851 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][7] ), 
        .B1(n6784), .B2(\IBusCachedPlugin_cache/banks_0[11][7] ), .ZN(n6746)
         );
  aoi22d1 U6852 ( .A1(n6754), .A2(\IBusCachedPlugin_cache/banks_0[3][7] ), 
        .B1(n6637), .B2(\IBusCachedPlugin_cache/banks_0[5][7] ), .ZN(n6745) );
  oai21d1 U6853 ( .B1(n6750), .B2(n6749), .A(n2356), .ZN(n6751) );
  oai21d1 U6854 ( .B1(n6800), .B2(n6752), .A(n6751), .ZN(n3985) );
  aoim22d1 U6855 ( .A1(n6753), .A2(n7113), .B1(n6997), .B2(
        memory_INSTRUCTION[7]), .Z(n3984) );
  aoi22d1 U6856 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][6] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][6] ), .ZN(n6758) );
  aoi22d1 U6857 ( .A1(n6790), .A2(\IBusCachedPlugin_cache/banks_0[12][6] ), 
        .B1(n6671), .B2(\IBusCachedPlugin_cache/banks_0[15][6] ), .ZN(n6757)
         );
  aoi22d1 U6858 ( .A1(n6772), .A2(\IBusCachedPlugin_cache/banks_0[2][6] ), 
        .B1(n6784), .B2(\IBusCachedPlugin_cache/banks_0[11][6] ), .ZN(n6756)
         );
  aoi22d1 U6859 ( .A1(n6754), .A2(\IBusCachedPlugin_cache/banks_0[3][6] ), 
        .B1(n6783), .B2(\IBusCachedPlugin_cache/banks_0[1][6] ), .ZN(n6755) );
  aoi22d1 U6860 ( .A1(n6537), .A2(\IBusCachedPlugin_cache/banks_0[14][6] ), 
        .B1(n6247), .B2(\IBusCachedPlugin_cache/banks_0[7][6] ), .ZN(n6762) );
  aoi22d1 U6861 ( .A1(n6791), .A2(\IBusCachedPlugin_cache/banks_0[5][6] ), 
        .B1(n7097), .B2(\IBusCachedPlugin_cache/banks_0[10][6] ), .ZN(n6761)
         );
  aoi22d1 U6862 ( .A1(n6628), .A2(\IBusCachedPlugin_cache/banks_0[6][6] ), 
        .B1(n6554), .B2(\IBusCachedPlugin_cache/banks_0[4][6] ), .ZN(n6760) );
  aoi22d1 U6863 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][6] ), 
        .B1(n7095), .B2(\IBusCachedPlugin_cache/banks_0[8][6] ), .ZN(n6759) );
  oai21d1 U6864 ( .B1(n6764), .B2(n6763), .A(n2356), .ZN(n6765) );
  oai21d1 U6865 ( .B1(n7107), .B2(n6766), .A(n6765), .ZN(n3983) );
  aoi22d1 U6866 ( .A1(n6652), .A2(\IBusCachedPlugin_cache/banks_0[11][5] ), 
        .B1(n6537), .B2(\IBusCachedPlugin_cache/banks_0[14][5] ), .ZN(n6771)
         );
  aoi22d1 U6867 ( .A1(n6767), .A2(\IBusCachedPlugin_cache/banks_0[1][5] ), 
        .B1(n6247), .B2(\IBusCachedPlugin_cache/banks_0[7][5] ), .ZN(n6770) );
  aoi22d1 U6868 ( .A1(n6628), .A2(\IBusCachedPlugin_cache/banks_0[6][5] ), 
        .B1(n7095), .B2(\IBusCachedPlugin_cache/banks_0[8][5] ), .ZN(n6769) );
  aoi22d1 U6869 ( .A1(n6637), .A2(\IBusCachedPlugin_cache/banks_0[5][5] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][5] ), .ZN(n6768) );
  aoi22d1 U6870 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][5] ), 
        .B1(n6671), .B2(\IBusCachedPlugin_cache/banks_0[15][5] ), .ZN(n6776)
         );
  aoi22d1 U6871 ( .A1(n6465), .A2(\IBusCachedPlugin_cache/banks_0[3][5] ), 
        .B1(n6554), .B2(\IBusCachedPlugin_cache/banks_0[4][5] ), .ZN(n6775) );
  aoi22d1 U6872 ( .A1(n6772), .A2(\IBusCachedPlugin_cache/banks_0[2][5] ), 
        .B1(n7097), .B2(\IBusCachedPlugin_cache/banks_0[10][5] ), .ZN(n6774)
         );
  aoi22d1 U6873 ( .A1(n6789), .A2(\IBusCachedPlugin_cache/banks_0[0][5] ), 
        .B1(n6790), .B2(\IBusCachedPlugin_cache/banks_0[12][5] ), .ZN(n6773)
         );
  oai21d1 U6874 ( .B1(n6778), .B2(n6777), .A(n2356), .ZN(n6779) );
  oai21d1 U6875 ( .B1(n6800), .B2(n6780), .A(n6779), .ZN(n3982) );
  aoi22d1 U6876 ( .A1(n6977), .A2(n6782), .B1(n6781), .B2(n6993), .ZN(n3980)
         );
  aoi22d1 U6877 ( .A1(n6465), .A2(\IBusCachedPlugin_cache/banks_0[3][4] ), 
        .B1(n6783), .B2(\IBusCachedPlugin_cache/banks_0[1][4] ), .ZN(n6788) );
  aoi22d1 U6878 ( .A1(n6772), .A2(\IBusCachedPlugin_cache/banks_0[2][4] ), 
        .B1(n6784), .B2(\IBusCachedPlugin_cache/banks_0[11][4] ), .ZN(n6787)
         );
  aoi22d1 U6879 ( .A1(n6672), .A2(\IBusCachedPlugin_cache/banks_0[13][4] ), 
        .B1(n6554), .B2(\IBusCachedPlugin_cache/banks_0[4][4] ), .ZN(n6786) );
  aoi22d1 U6880 ( .A1(n6537), .A2(\IBusCachedPlugin_cache/banks_0[14][4] ), 
        .B1(n6247), .B2(\IBusCachedPlugin_cache/banks_0[7][4] ), .ZN(n6785) );
  aoi22d1 U6881 ( .A1(n6789), .A2(\IBusCachedPlugin_cache/banks_0[0][4] ), 
        .B1(n7097), .B2(\IBusCachedPlugin_cache/banks_0[10][4] ), .ZN(n6795)
         );
  aoi22d1 U6882 ( .A1(n6791), .A2(\IBusCachedPlugin_cache/banks_0[5][4] ), 
        .B1(n6790), .B2(\IBusCachedPlugin_cache/banks_0[12][4] ), .ZN(n6794)
         );
  aoi22d1 U6883 ( .A1(n6651), .A2(\IBusCachedPlugin_cache/banks_0[9][4] ), 
        .B1(n6671), .B2(\IBusCachedPlugin_cache/banks_0[15][4] ), .ZN(n6793)
         );
  aoi22d1 U6884 ( .A1(n6628), .A2(\IBusCachedPlugin_cache/banks_0[6][4] ), 
        .B1(n7095), .B2(\IBusCachedPlugin_cache/banks_0[8][4] ), .ZN(n6792) );
  oai21d1 U6885 ( .B1(n6797), .B2(n6796), .A(n2356), .ZN(n6798) );
  oai21d1 U6886 ( .B1(n6800), .B2(n6799), .A(n6798), .ZN(n3979) );
  aoim22d1 U6887 ( .A1(n6801), .A2(n6926), .B1(n6996), .B2(memory_ENV_CTRL[0]), 
        .Z(n3978) );
  aoi22d1 U6888 ( .A1(n6889), .A2(n6803), .B1(n6802), .B2(n6997), .ZN(n3977)
         );
  aoim22d1 U6889 ( .A1(n6804), .A2(n7113), .B1(n6997), .B2(
        memory_REGFILE_WRITE_VALID), .Z(n3976) );
  aoim22d1 U6890 ( .A1(n6994), .A2(n7117), .B1(n6997), .B2(
        memory_MEMORY_ADDRESS_LOW[0]), .Z(n3975) );
  aoim22d1 U6891 ( .A1(n6981), .A2(n6997), .B1(n6997), .B2(
        memory_MEMORY_ADDRESS_LOW[1]), .Z(n3974) );
  nd02d0 U6892 ( .A1(execute_RS2[0]), .A2(n6972), .ZN(n6879) );
  oaim21d1 U6893 ( .B1(n7265), .B2(dBusWishbone_DAT_MOSI[0]), .A(n6879), .ZN(
        n3973) );
  inv0d1 U6894 ( .I(n6977), .ZN(n6965) );
  aoim22d1 U6895 ( .A1(n6805), .A2(n6972), .B1(n6965), .B2(
        dBusWishbone_ADR[29]), .Z(n3972) );
  aoim22d1 U6896 ( .A1(n6806), .A2(n6972), .B1(n6963), .B2(
        dBusWishbone_ADR[28]), .Z(n3971) );
  aoi22d1 U6897 ( .A1(n7085), .A2(n6808), .B1(n6807), .B2(n6862), .ZN(n3970)
         );
  aoi22d1 U6898 ( .A1(n6889), .A2(n6810), .B1(n6809), .B2(n6926), .ZN(n3969)
         );
  inv0d1 U6899 ( .I(n6977), .ZN(n6984) );
  aoim22d1 U6900 ( .A1(n6811), .A2(n6972), .B1(n6984), .B2(
        dBusWishbone_ADR[27]), .Z(n3968) );
  aoi22d1 U6901 ( .A1(n7090), .A2(n6813), .B1(n6812), .B2(n6862), .ZN(n3967)
         );
  aoi22d1 U6902 ( .A1(n7120), .A2(n6815), .B1(n6814), .B2(n7113), .ZN(n3966)
         );
  aoim22d1 U6903 ( .A1(n6816), .A2(n6972), .B1(n6984), .B2(
        dBusWishbone_ADR[26]), .Z(n3965) );
  aoi22d1 U6904 ( .A1(n7090), .A2(n6818), .B1(n6817), .B2(n6862), .ZN(n3964)
         );
  aoi22d1 U6905 ( .A1(n6889), .A2(n6820), .B1(n6819), .B2(n6926), .ZN(n3963)
         );
  aoim22d1 U6906 ( .A1(n6821), .A2(n6972), .B1(n6963), .B2(
        dBusWishbone_ADR[25]), .Z(n3962) );
  aoi22d1 U6907 ( .A1(n6939), .A2(n6823), .B1(n6822), .B2(n6862), .ZN(n3961)
         );
  aoi22d1 U6908 ( .A1(n6889), .A2(n6825), .B1(n6824), .B2(n6926), .ZN(n3960)
         );
  aoim22d1 U6909 ( .A1(n6826), .A2(n6972), .B1(n6965), .B2(
        dBusWishbone_ADR[24]), .Z(n3959) );
  aoi22d1 U6910 ( .A1(n7090), .A2(n6828), .B1(n6827), .B2(n6862), .ZN(n3958)
         );
  aoi22d1 U6911 ( .A1(n6889), .A2(n6830), .B1(n6829), .B2(n6926), .ZN(n3957)
         );
  aoim22d1 U6912 ( .A1(n6831), .A2(n6963), .B1(n6965), .B2(
        dBusWishbone_ADR[23]), .Z(n3956) );
  aoi22d1 U6913 ( .A1(n6939), .A2(n6833), .B1(n6832), .B2(n6862), .ZN(n3955)
         );
  aoi22d1 U6914 ( .A1(n6889), .A2(n6835), .B1(n6834), .B2(n6926), .ZN(n3954)
         );
  aoim22d1 U6915 ( .A1(n6836), .A2(n6963), .B1(n6984), .B2(
        dBusWishbone_ADR[22]), .Z(n3953) );
  aoi22d1 U6916 ( .A1(n7085), .A2(n6838), .B1(n6837), .B2(n6862), .ZN(n3952)
         );
  aoi22d1 U6917 ( .A1(n6889), .A2(n6840), .B1(n6839), .B2(n7113), .ZN(n3951)
         );
  aoim22d1 U6918 ( .A1(n6841), .A2(n6963), .B1(n6972), .B2(
        dBusWishbone_ADR[21]), .Z(n3950) );
  aoi22d1 U6919 ( .A1(n7090), .A2(n6843), .B1(n6842), .B2(n6862), .ZN(n3949)
         );
  aoi22d1 U6920 ( .A1(n6889), .A2(n6845), .B1(n6844), .B2(n6926), .ZN(n3948)
         );
  aoim22d1 U6921 ( .A1(n6846), .A2(n6963), .B1(n6963), .B2(
        dBusWishbone_ADR[20]), .Z(n3947) );
  aoi22d1 U6922 ( .A1(n6939), .A2(n6848), .B1(n6847), .B2(n6862), .ZN(n3946)
         );
  aoi22d1 U6923 ( .A1(n6889), .A2(n6850), .B1(n6849), .B2(n7113), .ZN(n3945)
         );
  aoim22d1 U6924 ( .A1(n6851), .A2(n6972), .B1(n6972), .B2(
        dBusWishbone_ADR[19]), .Z(n3944) );
  aoi22d1 U6925 ( .A1(n7090), .A2(n6853), .B1(n6852), .B2(n6862), .ZN(n3943)
         );
  aoi22d1 U6926 ( .A1(n6889), .A2(n6855), .B1(n6854), .B2(n6926), .ZN(n3942)
         );
  aoim22d1 U6927 ( .A1(n6856), .A2(n6963), .B1(n6963), .B2(
        dBusWishbone_ADR[18]), .Z(n3941) );
  aoi22d1 U6928 ( .A1(n6939), .A2(n6858), .B1(n6857), .B2(n6862), .ZN(n3940)
         );
  aoi22d1 U6929 ( .A1(n7120), .A2(n6860), .B1(n6859), .B2(n6926), .ZN(n3939)
         );
  aoim22d1 U6930 ( .A1(n6861), .A2(n6965), .B1(n6963), .B2(
        dBusWishbone_ADR[17]), .Z(n3938) );
  aoi22d1 U6931 ( .A1(n6939), .A2(n6864), .B1(n6863), .B2(n6862), .ZN(n3937)
         );
  aoi22d1 U6932 ( .A1(n6889), .A2(n6866), .B1(n6865), .B2(n6926), .ZN(n3936)
         );
  aoim22d1 U6933 ( .A1(n6867), .A2(n6965), .B1(n6920), .B2(
        dBusWishbone_ADR[16]), .Z(n3935) );
  aoi22d1 U6934 ( .A1(n6939), .A2(n6869), .B1(n6868), .B2(n6936), .ZN(n3934)
         );
  aoi22d1 U6935 ( .A1(n6889), .A2(n6871), .B1(n6870), .B2(n7113), .ZN(n3933)
         );
  aoim22d1 U6936 ( .A1(n6872), .A2(n6965), .B1(n6920), .B2(
        dBusWishbone_ADR[15]), .Z(n3932) );
  aoi22d1 U6937 ( .A1(n6939), .A2(n6874), .B1(n6873), .B2(n6936), .ZN(n3931)
         );
  aoi22d1 U6938 ( .A1(n7120), .A2(n6876), .B1(n6875), .B2(n6926), .ZN(n3930)
         );
  aoim22d1 U6939 ( .A1(n6877), .A2(n6965), .B1(n6984), .B2(
        dBusWishbone_ADR[14]), .Z(n3929) );
  aoi22d1 U6940 ( .A1(n6977), .A2(dBusWishbone_DAT_MOSI[16]), .B1(
        execute_RS2[16]), .B2(n6988), .ZN(n6878) );
  oai21d1 U6941 ( .B1(n6988), .B2(n6879), .A(n6878), .ZN(n3928) );
  aoi22d1 U6942 ( .A1(n7090), .A2(n6881), .B1(n6880), .B2(n6908), .ZN(n3927)
         );
  aoi22d1 U6943 ( .A1(n7120), .A2(n6883), .B1(n6882), .B2(n7113), .ZN(n3926)
         );
  aoim22d1 U6944 ( .A1(n6884), .A2(n6965), .B1(n6963), .B2(
        dBusWishbone_ADR[13]), .Z(n3925) );
  aoi22d1 U6945 ( .A1(n6939), .A2(n6886), .B1(n6885), .B2(n6936), .ZN(n3924)
         );
  aoi22d1 U6946 ( .A1(n6889), .A2(n6888), .B1(n6887), .B2(n7113), .ZN(n3923)
         );
  aoim22d1 U6947 ( .A1(n6890), .A2(n6965), .B1(n6963), .B2(
        dBusWishbone_ADR[12]), .Z(n3922) );
  aoi22d1 U6948 ( .A1(n6893), .A2(n6892), .B1(n6891), .B2(n6936), .ZN(n3921)
         );
  aoi22d1 U6949 ( .A1(n7120), .A2(n6895), .B1(n6894), .B2(n6926), .ZN(n3920)
         );
  aoim22d1 U6950 ( .A1(n6896), .A2(n6984), .B1(n6972), .B2(
        dBusWishbone_ADR[11]), .Z(n3919) );
  aoim22d1 U6951 ( .A1(n6897), .A2(n6965), .B1(n6965), .B2(
        dBusWishbone_ADR[10]), .Z(n3918) );
  aoi22d1 U6952 ( .A1(n6939), .A2(n6899), .B1(n6898), .B2(n6908), .ZN(n3917)
         );
  aoi22d1 U6953 ( .A1(n7120), .A2(n6901), .B1(n6900), .B2(n7113), .ZN(n3916)
         );
  aoim22d1 U6954 ( .A1(n6902), .A2(n6984), .B1(n6984), .B2(dBusWishbone_ADR[9]), .Z(n3915) );
  aoi22d1 U6955 ( .A1(n7090), .A2(n6904), .B1(n6903), .B2(n6908), .ZN(n3914)
         );
  aoi22d1 U6956 ( .A1(n7120), .A2(n6906), .B1(n6905), .B2(n7113), .ZN(n3913)
         );
  aoim22d1 U6957 ( .A1(n6907), .A2(n6963), .B1(n6972), .B2(dBusWishbone_ADR[8]), .Z(n3912) );
  aoi22d1 U6958 ( .A1(n6939), .A2(n6910), .B1(n6909), .B2(n6908), .ZN(n3911)
         );
  aoi22d1 U6959 ( .A1(n7120), .A2(n6912), .B1(n6911), .B2(n6926), .ZN(n3910)
         );
  aoim22d1 U6960 ( .A1(n6913), .A2(n6984), .B1(n6965), .B2(dBusWishbone_ADR[7]), .Z(n3909) );
  aoi22d1 U6961 ( .A1(n6939), .A2(n6915), .B1(n6914), .B2(n6936), .ZN(n3908)
         );
  aoi22d1 U6962 ( .A1(n7120), .A2(n6917), .B1(n6916), .B2(n7113), .ZN(n3907)
         );
  aoim22d1 U6963 ( .A1(n6918), .A2(n6984), .B1(n6972), .B2(dBusWishbone_ADR[6]), .Z(n3906) );
  nd03d0 U6964 ( .A1(execute_ALU_BITWISE_CTRL[1]), .A2(n6920), .A3(n6919), 
        .ZN(n6992) );
  inv0d0 U6965 ( .I(execute_RS2[8]), .ZN(n6923) );
  aoi22d1 U6966 ( .A1(n6977), .A2(dBusWishbone_DAT_MOSI[24]), .B1(
        execute_RS2[24]), .B2(n6988), .ZN(n6922) );
  oai211d1 U6967 ( .C1(n6992), .C2(n6923), .A(n6922), .B(n6921), .ZN(n3904) );
  aoi22d1 U6968 ( .A1(n7085), .A2(n6925), .B1(n6924), .B2(n6936), .ZN(n3903)
         );
  aoi22d1 U6969 ( .A1(n7120), .A2(n6928), .B1(n6927), .B2(n6926), .ZN(n3902)
         );
  aoim22d1 U6970 ( .A1(n6929), .A2(n6965), .B1(n6963), .B2(dBusWishbone_ADR[5]), .Z(n3901) );
  nd02d0 U6971 ( .A1(execute_RS2[7]), .A2(n6965), .ZN(n6931) );
  oaim21d1 U6972 ( .B1(n7265), .B2(dBusWishbone_DAT_MOSI[7]), .A(n6931), .ZN(
        n3900) );
  inv0d0 U6973 ( .I(execute_RS2[23]), .ZN(n6932) );
  inv0d0 U6974 ( .I(dBusWishbone_DAT_MOSI[23]), .ZN(n6930) );
  oai222d1 U6975 ( .A1(n6932), .A2(n6986), .B1(n6931), .B2(
        _zz__zz_execute_BranchPlugin_branch_src2[12]), .C1(n6984), .C2(n6930), 
        .ZN(n3898) );
  inv0d0 U6976 ( .I(execute_RS2[15]), .ZN(n6935) );
  aoi22d1 U6977 ( .A1(n6977), .A2(dBusWishbone_DAT_MOSI[31]), .B1(
        execute_RS2[31]), .B2(n6988), .ZN(n6934) );
  oai211d1 U6978 ( .C1(n6992), .C2(n6935), .A(n6934), .B(n6933), .ZN(n3897) );
  aoi22d1 U6979 ( .A1(n6939), .A2(n6938), .B1(n6937), .B2(n6936), .ZN(n3896)
         );
  aoi22d1 U6980 ( .A1(n7004), .A2(n6941), .B1(n6940), .B2(n7113), .ZN(n3895)
         );
  aoim22d1 U6981 ( .A1(n6943), .A2(n6965), .B1(n6963), .B2(dBusWishbone_ADR[4]), .Z(n3894) );
  nd02d0 U6982 ( .A1(execute_RS2[6]), .A2(n6965), .ZN(n6945) );
  oaim21d1 U6983 ( .B1(n7265), .B2(dBusWishbone_DAT_MOSI[6]), .A(n6945), .ZN(
        n3893) );
  aoi22d1 U6984 ( .A1(n7265), .A2(dBusWishbone_DAT_MOSI[22]), .B1(
        execute_RS2[22]), .B2(n6988), .ZN(n6944) );
  oai21d1 U6985 ( .B1(n6988), .B2(n6945), .A(n6944), .ZN(n3891) );
  inv0d0 U6986 ( .I(execute_RS2[14]), .ZN(n6948) );
  aoi22d1 U6987 ( .A1(dBusWishbone_CYC), .A2(dBusWishbone_DAT_MOSI[30]), .B1(
        execute_RS2[30]), .B2(n6988), .ZN(n6947) );
  oai211d1 U6988 ( .C1(n6992), .C2(n6948), .A(n6947), .B(n6946), .ZN(n3890) );
  aoim22d1 U6989 ( .A1(n6949), .A2(n6963), .B1(n6993), .B2(dBusWishbone_ADR[3]), .Z(n3889) );
  nd02d0 U6990 ( .A1(execute_RS2[5]), .A2(n6963), .ZN(n6951) );
  oaim21d1 U6991 ( .B1(n7265), .B2(dBusWishbone_DAT_MOSI[5]), .A(n6951), .ZN(
        n3888) );
  inv0d0 U6992 ( .I(execute_RS2[21]), .ZN(n6952) );
  inv0d0 U6993 ( .I(dBusWishbone_DAT_MOSI[21]), .ZN(n6950) );
  oai222d1 U6994 ( .A1(n6952), .A2(n6986), .B1(n6951), .B2(
        _zz__zz_execute_BranchPlugin_branch_src2[12]), .C1(n6984), .C2(n6950), 
        .ZN(n3886) );
  inv0d0 U6995 ( .I(execute_RS2[13]), .ZN(n6955) );
  aoi22d1 U6996 ( .A1(dBusWishbone_CYC), .A2(dBusWishbone_DAT_MOSI[29]), .B1(
        execute_RS2[29]), .B2(n6988), .ZN(n6954) );
  oai211d1 U6997 ( .C1(n6992), .C2(n6955), .A(n6954), .B(n6953), .ZN(n3885) );
  aoim22d1 U6998 ( .A1(n6956), .A2(n6963), .B1(n6993), .B2(dBusWishbone_ADR[2]), .Z(n3884) );
  nd02d0 U6999 ( .A1(execute_RS2[4]), .A2(n6972), .ZN(n6958) );
  oaim21d1 U7000 ( .B1(n7265), .B2(dBusWishbone_DAT_MOSI[4]), .A(n6958), .ZN(
        n3883) );
  inv0d0 U7001 ( .I(execute_RS2[20]), .ZN(n6959) );
  inv0d0 U7002 ( .I(dBusWishbone_DAT_MOSI[20]), .ZN(n6957) );
  oai222d1 U7003 ( .A1(n6959), .A2(n6986), .B1(n6958), .B2(
        _zz__zz_execute_BranchPlugin_branch_src2[12]), .C1(n6984), .C2(n6957), 
        .ZN(n3881) );
  inv0d0 U7004 ( .I(execute_RS2[12]), .ZN(n6962) );
  aoi22d1 U7005 ( .A1(dBusWishbone_CYC), .A2(dBusWishbone_DAT_MOSI[28]), .B1(
        execute_RS2[28]), .B2(n6988), .ZN(n6961) );
  oai211d1 U7006 ( .C1(n6992), .C2(n6962), .A(n6961), .B(n6960), .ZN(n3880) );
  aoim22d1 U7007 ( .A1(n6964), .A2(n6963), .B1(n6993), .B2(dBusWishbone_ADR[1]), .Z(n3879) );
  nd02d0 U7008 ( .A1(execute_RS2[3]), .A2(n6965), .ZN(n6967) );
  oaim21d1 U7009 ( .B1(n7265), .B2(dBusWishbone_DAT_MOSI[3]), .A(n6967), .ZN(
        n3878) );
  inv0d0 U7010 ( .I(execute_RS2[19]), .ZN(n6968) );
  inv0d0 U7011 ( .I(dBusWishbone_DAT_MOSI[19]), .ZN(n6966) );
  oai222d1 U7012 ( .A1(n6968), .A2(n6986), .B1(n6967), .B2(
        _zz__zz_execute_BranchPlugin_branch_src2[12]), .C1(n6984), .C2(n6966), 
        .ZN(n3876) );
  inv0d0 U7013 ( .I(execute_RS2[11]), .ZN(n6971) );
  aoi22d1 U7014 ( .A1(dBusWishbone_CYC), .A2(dBusWishbone_DAT_MOSI[27]), .B1(
        execute_RS2[27]), .B2(n6988), .ZN(n6970) );
  oai211d1 U7015 ( .C1(n6992), .C2(n6971), .A(n6970), .B(n6969), .ZN(n3875) );
  aoim22d1 U7016 ( .A1(n6973), .A2(n6972), .B1(n6993), .B2(dBusWishbone_ADR[0]), .Z(n3874) );
  nd02d0 U7017 ( .A1(execute_RS2[2]), .A2(n6984), .ZN(n6975) );
  oaim21d1 U7018 ( .B1(n7265), .B2(dBusWishbone_DAT_MOSI[2]), .A(n6975), .ZN(
        n3873) );
  inv0d0 U7019 ( .I(execute_RS2[18]), .ZN(n6976) );
  inv0d0 U7020 ( .I(dBusWishbone_DAT_MOSI[18]), .ZN(n6974) );
  oai222d1 U7021 ( .A1(n6976), .A2(n6986), .B1(n6975), .B2(
        _zz__zz_execute_BranchPlugin_branch_src2[12]), .C1(n6984), .C2(n6974), 
        .ZN(n3871) );
  inv0d0 U7022 ( .I(execute_RS2[10]), .ZN(n6980) );
  aoi22d1 U7023 ( .A1(n6977), .A2(dBusWishbone_DAT_MOSI[26]), .B1(
        execute_RS2[26]), .B2(n6988), .ZN(n6979) );
  oai211d1 U7024 ( .C1(n6992), .C2(n6980), .A(n6979), .B(n6978), .ZN(n3870) );
  aoi22d1 U7025 ( .A1(dBusWishbone_CYC), .A2(n6982), .B1(n6981), .B2(n6993), 
        .ZN(n3869) );
  nd02d0 U7026 ( .A1(execute_RS2[1]), .A2(n6984), .ZN(n6985) );
  oaim21d1 U7027 ( .B1(n7265), .B2(dBusWishbone_DAT_MOSI[1]), .A(n6985), .ZN(
        n3868) );
  inv0d0 U7028 ( .I(execute_RS2[17]), .ZN(n6987) );
  inv0d0 U7029 ( .I(dBusWishbone_DAT_MOSI[17]), .ZN(n6983) );
  oai222d1 U7030 ( .A1(n6987), .A2(n6986), .B1(n6985), .B2(
        _zz__zz_execute_BranchPlugin_branch_src2[12]), .C1(n6984), .C2(n6983), 
        .ZN(n3866) );
  inv0d0 U7031 ( .I(execute_RS2[9]), .ZN(n6991) );
  aoi22d1 U7032 ( .A1(dBusWishbone_CYC), .A2(dBusWishbone_DAT_MOSI[25]), .B1(
        execute_RS2[25]), .B2(n6988), .ZN(n6990) );
  oai211d1 U7033 ( .C1(n6992), .C2(n6991), .A(n6990), .B(n6989), .ZN(n3865) );
  aoi22d1 U7034 ( .A1(dBusWishbone_CYC), .A2(n6995), .B1(n6994), .B2(n6993), 
        .ZN(n3864) );
  aoim22d1 U7035 ( .A1(n6998), .A2(n6997), .B1(n6996), .B2(
        memory_ALIGNEMENT_FAULT), .Z(n3863) );
  aoi22d1 U7036 ( .A1(n7085), .A2(n7001), .B1(n7000), .B2(n6999), .ZN(n3862)
         );
  aoi22d1 U7037 ( .A1(n7004), .A2(n7003), .B1(n7002), .B2(n7113), .ZN(n3861)
         );
  nd02d1 U7038 ( .A1(n7007), .A2(n7005), .ZN(n7087) );
  inv0d0 U7039 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[0] ), .ZN(
        n7009) );
  oai222d1 U7040 ( .A1(n7010), .A2(n7087), .B1(n7009), .B2(n7107), .C1(n7077), 
        .C2(n7008), .ZN(n3860) );
  buffd1 U7041 ( .I(n7087), .Z(n7092) );
  oai222d1 U7042 ( .A1(n7013), .A2(n7077), .B1(n7012), .B2(n7085), .C1(n7011), 
        .C2(n7092), .ZN(n3859) );
  oai222d1 U7043 ( .A1(n7016), .A2(n7077), .B1(n7015), .B2(n7085), .C1(n7014), 
        .C2(n7092), .ZN(n3858) );
  oai222d1 U7044 ( .A1(n7019), .A2(n7092), .B1(n7018), .B2(n6800), .C1(n7017), 
        .C2(n7077), .ZN(n3857) );
  oai222d1 U7045 ( .A1(n7022), .A2(n7092), .B1(n7021), .B2(n7090), .C1(n7020), 
        .C2(n7077), .ZN(n3856) );
  oai222d1 U7046 ( .A1(n7025), .A2(n7077), .B1(n7024), .B2(n7085), .C1(n7023), 
        .C2(n7092), .ZN(n3855) );
  oai222d1 U7047 ( .A1(n7028), .A2(n7092), .B1(n7027), .B2(n7107), .C1(n7026), 
        .C2(n7077), .ZN(n3854) );
  inv0d0 U7048 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[21] ), .ZN(
        n7030) );
  oai222d1 U7049 ( .A1(n7031), .A2(n7087), .B1(n7030), .B2(n7085), .C1(n7029), 
        .C2(n7077), .ZN(n3853) );
  oai222d1 U7050 ( .A1(n7034), .A2(n7087), .B1(n7033), .B2(n7090), .C1(n7032), 
        .C2(n7077), .ZN(n3852) );
  oai222d1 U7051 ( .A1(n7037), .A2(n7077), .B1(n7036), .B2(n2356), .C1(n7035), 
        .C2(n7092), .ZN(n3851) );
  oai222d1 U7052 ( .A1(n7040), .A2(n7092), .B1(n7039), .B2(n7107), .C1(n7038), 
        .C2(n7077), .ZN(n3850) );
  oai222d1 U7053 ( .A1(n7043), .A2(n7092), .B1(n7042), .B2(n7085), .C1(n7041), 
        .C2(n7077), .ZN(n3849) );
  inv0d0 U7054 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[16] ), .ZN(
        n7045) );
  oai222d1 U7055 ( .A1(n7046), .A2(n7087), .B1(n7045), .B2(n7085), .C1(n7044), 
        .C2(n7077), .ZN(n3848) );
  oai222d1 U7056 ( .A1(n7049), .A2(n7077), .B1(n7048), .B2(n6800), .C1(n7047), 
        .C2(n7092), .ZN(n3847) );
  oai222d1 U7057 ( .A1(n7052), .A2(n7092), .B1(n7051), .B2(n7107), .C1(n7050), 
        .C2(n7077), .ZN(n3846) );
  inv0d0 U7058 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[13] ), .ZN(
        n7054) );
  oai222d1 U7059 ( .A1(n7055), .A2(n7077), .B1(n7054), .B2(n7085), .C1(n7053), 
        .C2(n7087), .ZN(n3845) );
  inv0d0 U7060 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[12] ), .ZN(
        n7057) );
  oai222d1 U7061 ( .A1(n7058), .A2(n7077), .B1(n7057), .B2(n2356), .C1(n7056), 
        .C2(n7092), .ZN(n3844) );
  oai222d1 U7062 ( .A1(n7061), .A2(n7077), .B1(n7060), .B2(n7090), .C1(n7059), 
        .C2(n7087), .ZN(n3843) );
  oai222d1 U7063 ( .A1(n7064), .A2(n7087), .B1(n7063), .B2(n7090), .C1(n7062), 
        .C2(n7077), .ZN(n3842) );
  inv0d0 U7064 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[9] ), .ZN(
        n7066) );
  oai222d1 U7065 ( .A1(n7067), .A2(n7077), .B1(n7066), .B2(n6939), .C1(n7065), 
        .C2(n7092), .ZN(n3841) );
  oai222d1 U7066 ( .A1(n7070), .A2(n7077), .B1(n7069), .B2(n7090), .C1(n7068), 
        .C2(n7092), .ZN(n3840) );
  oai222d1 U7067 ( .A1(n7073), .A2(n7077), .B1(n7072), .B2(n7090), .C1(n7071), 
        .C2(n7092), .ZN(n3839) );
  inv0d0 U7068 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[6] ), .ZN(
        n7075) );
  oai222d1 U7069 ( .A1(n7076), .A2(n7092), .B1(n7075), .B2(n7085), .C1(n7074), 
        .C2(n7077), .ZN(n3838) );
  oai222d1 U7070 ( .A1(n7080), .A2(n7087), .B1(n7079), .B2(n7090), .C1(n7078), 
        .C2(n7077), .ZN(n3837) );
  inv0d0 U7071 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[4] ), .ZN(
        n7082) );
  oai222d1 U7072 ( .A1(n7083), .A2(n7087), .B1(n7082), .B2(n7085), .C1(n7081), 
        .C2(n7077), .ZN(n3836) );
  inv0d0 U7073 ( .I(\IBusCachedPlugin_cache/_zz_ways_0_tags_port1[3] ), .ZN(
        n7086) );
  oai222d1 U7074 ( .A1(n7088), .A2(n7087), .B1(n7086), .B2(n7085), .C1(n7084), 
        .C2(n7077), .ZN(n3835) );
  oai222d1 U7075 ( .A1(n7093), .A2(n7092), .B1(n7091), .B2(n7090), .C1(n7089), 
        .C2(n7077), .ZN(n3834) );
  aoi22d1 U7076 ( .A1(n7094), .A2(\IBusCachedPlugin_cache/banks_0[0][1] ), 
        .B1(n6651), .B2(\IBusCachedPlugin_cache/banks_0[9][1] ), .ZN(n7101) );
  aoi22d1 U7077 ( .A1(n6628), .A2(\IBusCachedPlugin_cache/banks_0[6][1] ), 
        .B1(n7095), .B2(\IBusCachedPlugin_cache/banks_0[8][1] ), .ZN(n7100) );
  aoi22d1 U7078 ( .A1(n7096), .A2(\IBusCachedPlugin_cache/banks_0[2][1] ), 
        .B1(n6475), .B2(\IBusCachedPlugin_cache/banks_0[12][1] ), .ZN(n7099)
         );
  aoi22d1 U7079 ( .A1(n7097), .A2(\IBusCachedPlugin_cache/banks_0[10][1] ), 
        .B1(n6671), .B2(\IBusCachedPlugin_cache/banks_0[15][1] ), .ZN(n7098)
         );
  aoi22d1 U7080 ( .A1(n6637), .A2(\IBusCachedPlugin_cache/banks_0[5][1] ), 
        .B1(n6672), .B2(\IBusCachedPlugin_cache/banks_0[13][1] ), .ZN(n7106)
         );
  aoi22d1 U7081 ( .A1(n6652), .A2(\IBusCachedPlugin_cache/banks_0[11][1] ), 
        .B1(n6247), .B2(\IBusCachedPlugin_cache/banks_0[7][1] ), .ZN(n7105) );
  aoi22d1 U7082 ( .A1(n6767), .A2(\IBusCachedPlugin_cache/banks_0[1][1] ), 
        .B1(n7102), .B2(\IBusCachedPlugin_cache/banks_0[4][1] ), .ZN(n7104) );
  aoi22d1 U7083 ( .A1(n6465), .A2(\IBusCachedPlugin_cache/banks_0[3][1] ), 
        .B1(n6537), .B2(\IBusCachedPlugin_cache/banks_0[14][1] ), .ZN(n7103)
         );
  oai21d1 U7084 ( .B1(n7109), .B2(n7108), .A(n7107), .ZN(n7110) );
  oai21d1 U7085 ( .B1(n7112), .B2(n7111), .A(n7110), .ZN(n3833) );
  aoi22d1 U7086 ( .A1(n7116), .A2(n7115), .B1(n7114), .B2(n7113), .ZN(n3832)
         );
  aoi22d1 U7087 ( .A1(n7120), .A2(n7119), .B1(n7118), .B2(n7117), .ZN(n3831)
         );
endmodule


