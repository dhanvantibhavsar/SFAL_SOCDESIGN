module housekeeping ( VPWR, VGND, wb_clk_i, wb_adr_i, wb_dat_i, wb_sel_i, 
        wb_we_i, wb_cyc_i, wb_stb_i, wb_ack_o, wb_dat_o, porb, pll_ena, 
        pll_dco_ena, pll_div, pll_sel, pll90_sel, pll_trim, pll_bypass, 
        qspi_enabled, uart_enabled, spi_enabled, debug_mode, ser_tx, ser_rx, 
        spi_sdi, spi_csb, spi_sck, spi_sdo, spi_sdoenb, irq, reset, 
        serial_clock, serial_load, serial_resetn, serial_data_1, serial_data_2, 
        mgmt_gpio_in, mgmt_gpio_out, mgmt_gpio_oeb, pwr_ctrl_out, trap, 
        user_clock, mask_rev_in, spimemio_flash_csb, spimemio_flash_clk, 
        spimemio_flash_io0_oeb, spimemio_flash_io1_oeb, spimemio_flash_io2_oeb, 
        spimemio_flash_io3_oeb, spimemio_flash_io0_do, spimemio_flash_io1_do, 
        spimemio_flash_io2_do, spimemio_flash_io3_do, spimemio_flash_io0_di, 
        spimemio_flash_io1_di, spimemio_flash_io2_di, spimemio_flash_io3_di, 
        debug_in, debug_out, debug_oeb, pad_flash_csb, pad_flash_csb_oeb, 
        pad_flash_clk, pad_flash_clk_oeb, pad_flash_io0_oeb, pad_flash_io1_oeb, 
        pad_flash_io0_ieb, pad_flash_io1_ieb, pad_flash_io0_do, 
        pad_flash_io1_do, pad_flash_io0_di, pad_flash_io1_di, usr1_vcc_pwrgood, 
        usr2_vcc_pwrgood, usr1_vdd_pwrgood, usr2_vdd_pwrgood, wb_rstn_i_BAR );
  input [31:0] wb_adr_i;
  input [31:0] wb_dat_i;
  input [3:0] wb_sel_i;
  output [31:0] wb_dat_o;
  output [4:0] pll_div;
  output [2:0] pll_sel;
  output [2:0] pll90_sel;
  output [25:0] pll_trim;
  output [2:0] irq;
  input [37:0] mgmt_gpio_in;
  output [37:0] mgmt_gpio_out;
  output [37:0] mgmt_gpio_oeb;
  output [3:0] pwr_ctrl_out;
  input [31:0] mask_rev_in;
  input wb_clk_i, wb_we_i, wb_cyc_i, wb_stb_i, porb, qspi_enabled,
         uart_enabled, spi_enabled, debug_mode, ser_tx, spi_csb, spi_sck,
         spi_sdo, spi_sdoenb, trap, user_clock, spimemio_flash_csb,
         spimemio_flash_clk, spimemio_flash_io0_oeb, spimemio_flash_io1_oeb,
         spimemio_flash_io2_oeb, spimemio_flash_io3_oeb, spimemio_flash_io0_do,
         spimemio_flash_io1_do, spimemio_flash_io2_do, spimemio_flash_io3_do,
         debug_out, debug_oeb, pad_flash_io0_di, pad_flash_io1_di,
         usr1_vcc_pwrgood, usr2_vcc_pwrgood, usr1_vdd_pwrgood,
         usr2_vdd_pwrgood, wb_rstn_i_BAR;
  output wb_ack_o, pll_ena, pll_dco_ena, pll_bypass, ser_rx, spi_sdi, reset,
         serial_clock, serial_load, serial_resetn, serial_data_1,
         serial_data_2, spimemio_flash_io0_di, spimemio_flash_io1_di,
         spimemio_flash_io2_di, spimemio_flash_io3_di, debug_in, pad_flash_csb,
         pad_flash_csb_oeb, pad_flash_clk, pad_flash_clk_oeb,
         pad_flash_io0_oeb, pad_flash_io1_oeb, pad_flash_io0_ieb,
         pad_flash_io1_ieb, pad_flash_io0_do, pad_flash_io1_do;
  inout VPWR,  VGND;
  wire   wb_rstn_i, n429, n430, n431, n432, n3390, reset_reg,
         pass_thru_mgmt_delay, pass_thru_mgmt, \gpio_configure[37][12] ,
         \gpio_configure[37][11] , \gpio_configure[37][10] ,
         \gpio_configure[37][9] , \gpio_configure[37][8] ,
         \gpio_configure[37][7] , \gpio_configure[37][6] ,
         \gpio_configure[37][5] , \gpio_configure[37][4] ,
         \gpio_configure[37][3] , \gpio_configure[37][2] ,
         \gpio_configure[37][1] , \gpio_configure[37][0] ,
         \gpio_configure[36][12] , \gpio_configure[36][11] ,
         \gpio_configure[36][10] , \gpio_configure[36][9] ,
         \gpio_configure[36][8] , \gpio_configure[36][7] ,
         \gpio_configure[36][6] , \gpio_configure[36][5] ,
         \gpio_configure[36][4] , \gpio_configure[36][3] ,
         \gpio_configure[36][2] , \gpio_configure[36][1] ,
         \gpio_configure[36][0] , \gpio_configure[35][12] ,
         \gpio_configure[35][11] , \gpio_configure[35][10] ,
         \gpio_configure[35][9] , \gpio_configure[35][8] ,
         \gpio_configure[35][7] , \gpio_configure[35][6] ,
         \gpio_configure[35][5] , \gpio_configure[35][4] ,
         \gpio_configure[35][3] , \gpio_configure[35][2] ,
         \gpio_configure[35][1] , \gpio_configure[35][0] ,
         \gpio_configure[34][12] , \gpio_configure[34][11] ,
         \gpio_configure[34][10] , \gpio_configure[34][9] ,
         \gpio_configure[34][8] , \gpio_configure[34][7] ,
         \gpio_configure[34][6] , \gpio_configure[34][5] ,
         \gpio_configure[34][4] , \gpio_configure[34][3] ,
         \gpio_configure[34][2] , \gpio_configure[34][1] ,
         \gpio_configure[34][0] , \gpio_configure[33][12] ,
         \gpio_configure[33][11] , \gpio_configure[33][10] ,
         \gpio_configure[33][9] , \gpio_configure[33][8] ,
         \gpio_configure[33][7] , \gpio_configure[33][6] ,
         \gpio_configure[33][5] , \gpio_configure[33][4] ,
         \gpio_configure[33][3] , \gpio_configure[33][2] ,
         \gpio_configure[33][1] , \gpio_configure[33][0] ,
         \gpio_configure[32][12] , \gpio_configure[32][11] ,
         \gpio_configure[32][10] , \gpio_configure[32][9] ,
         \gpio_configure[32][8] , \gpio_configure[32][7] ,
         \gpio_configure[32][6] , \gpio_configure[32][5] ,
         \gpio_configure[32][4] , \gpio_configure[32][3] ,
         \gpio_configure[32][2] , \gpio_configure[32][1] ,
         \gpio_configure[32][0] , \gpio_configure[31][12] ,
         \gpio_configure[31][11] , \gpio_configure[31][10] ,
         \gpio_configure[31][9] , \gpio_configure[31][8] ,
         \gpio_configure[31][7] , \gpio_configure[31][6] ,
         \gpio_configure[31][5] , \gpio_configure[31][4] ,
         \gpio_configure[31][3] , \gpio_configure[31][2] ,
         \gpio_configure[31][1] , \gpio_configure[31][0] ,
         \gpio_configure[30][12] , \gpio_configure[30][11] ,
         \gpio_configure[30][10] , \gpio_configure[30][9] ,
         \gpio_configure[30][8] , \gpio_configure[30][7] ,
         \gpio_configure[30][6] , \gpio_configure[30][5] ,
         \gpio_configure[30][4] , \gpio_configure[30][3] ,
         \gpio_configure[30][2] , \gpio_configure[30][1] ,
         \gpio_configure[30][0] , \gpio_configure[29][12] ,
         \gpio_configure[29][11] , \gpio_configure[29][10] ,
         \gpio_configure[29][9] , \gpio_configure[29][8] ,
         \gpio_configure[29][7] , \gpio_configure[29][6] ,
         \gpio_configure[29][5] , \gpio_configure[29][4] ,
         \gpio_configure[29][3] , \gpio_configure[29][2] ,
         \gpio_configure[29][1] , \gpio_configure[29][0] ,
         \gpio_configure[28][12] , \gpio_configure[28][11] ,
         \gpio_configure[28][10] , \gpio_configure[28][9] ,
         \gpio_configure[28][8] , \gpio_configure[28][7] ,
         \gpio_configure[28][6] , \gpio_configure[28][5] ,
         \gpio_configure[28][4] , \gpio_configure[28][3] ,
         \gpio_configure[28][2] , \gpio_configure[28][1] ,
         \gpio_configure[28][0] , \gpio_configure[27][12] ,
         \gpio_configure[27][11] , \gpio_configure[27][10] ,
         \gpio_configure[27][9] , \gpio_configure[27][8] ,
         \gpio_configure[27][7] , \gpio_configure[27][6] ,
         \gpio_configure[27][5] , \gpio_configure[27][4] ,
         \gpio_configure[27][3] , \gpio_configure[27][2] ,
         \gpio_configure[27][1] , \gpio_configure[27][0] ,
         \gpio_configure[26][12] , \gpio_configure[26][11] ,
         \gpio_configure[26][10] , \gpio_configure[26][9] ,
         \gpio_configure[26][8] , \gpio_configure[26][7] ,
         \gpio_configure[26][6] , \gpio_configure[26][5] ,
         \gpio_configure[26][4] , \gpio_configure[26][3] ,
         \gpio_configure[26][2] , \gpio_configure[26][1] ,
         \gpio_configure[26][0] , \gpio_configure[25][12] ,
         \gpio_configure[25][11] , \gpio_configure[25][10] ,
         \gpio_configure[25][9] , \gpio_configure[25][8] ,
         \gpio_configure[25][7] , \gpio_configure[25][6] ,
         \gpio_configure[25][5] , \gpio_configure[25][4] ,
         \gpio_configure[25][3] , \gpio_configure[25][2] ,
         \gpio_configure[25][1] , \gpio_configure[25][0] ,
         \gpio_configure[24][12] , \gpio_configure[24][11] ,
         \gpio_configure[24][10] , \gpio_configure[24][9] ,
         \gpio_configure[24][8] , \gpio_configure[24][7] ,
         \gpio_configure[24][6] , \gpio_configure[24][5] ,
         \gpio_configure[24][4] , \gpio_configure[24][3] ,
         \gpio_configure[24][2] , \gpio_configure[24][1] ,
         \gpio_configure[24][0] , \gpio_configure[23][12] ,
         \gpio_configure[23][11] , \gpio_configure[23][10] ,
         \gpio_configure[23][9] , \gpio_configure[23][8] ,
         \gpio_configure[23][7] , \gpio_configure[23][6] ,
         \gpio_configure[23][5] , \gpio_configure[23][4] ,
         \gpio_configure[23][3] , \gpio_configure[23][2] ,
         \gpio_configure[23][1] , \gpio_configure[23][0] ,
         \gpio_configure[22][12] , \gpio_configure[22][11] ,
         \gpio_configure[22][10] , \gpio_configure[22][9] ,
         \gpio_configure[22][8] , \gpio_configure[22][7] ,
         \gpio_configure[22][6] , \gpio_configure[22][5] ,
         \gpio_configure[22][4] , \gpio_configure[22][3] ,
         \gpio_configure[22][2] , \gpio_configure[22][1] ,
         \gpio_configure[22][0] , \gpio_configure[21][12] ,
         \gpio_configure[21][11] , \gpio_configure[21][10] ,
         \gpio_configure[21][9] , \gpio_configure[21][8] ,
         \gpio_configure[21][7] , \gpio_configure[21][6] ,
         \gpio_configure[21][5] , \gpio_configure[21][4] ,
         \gpio_configure[21][3] , \gpio_configure[21][2] ,
         \gpio_configure[21][1] , \gpio_configure[21][0] ,
         \gpio_configure[20][12] , \gpio_configure[20][11] ,
         \gpio_configure[20][10] , \gpio_configure[20][9] ,
         \gpio_configure[20][8] , \gpio_configure[20][7] ,
         \gpio_configure[20][6] , \gpio_configure[20][5] ,
         \gpio_configure[20][4] , \gpio_configure[20][3] ,
         \gpio_configure[20][2] , \gpio_configure[20][1] ,
         \gpio_configure[20][0] , \gpio_configure[19][12] ,
         \gpio_configure[19][11] , \gpio_configure[19][10] ,
         \gpio_configure[19][9] , \gpio_configure[19][8] ,
         \gpio_configure[19][7] , \gpio_configure[19][6] ,
         \gpio_configure[19][5] , \gpio_configure[19][4] ,
         \gpio_configure[19][3] , \gpio_configure[19][2] ,
         \gpio_configure[19][1] , \gpio_configure[19][0] ,
         \gpio_configure[18][12] , \gpio_configure[18][11] ,
         \gpio_configure[18][10] , \gpio_configure[18][9] ,
         \gpio_configure[18][8] , \gpio_configure[18][7] ,
         \gpio_configure[18][6] , \gpio_configure[18][5] ,
         \gpio_configure[18][4] , \gpio_configure[18][3] ,
         \gpio_configure[18][2] , \gpio_configure[18][1] ,
         \gpio_configure[18][0] , \gpio_configure[17][12] ,
         \gpio_configure[17][11] , \gpio_configure[17][10] ,
         \gpio_configure[17][9] , \gpio_configure[17][8] ,
         \gpio_configure[17][7] , \gpio_configure[17][6] ,
         \gpio_configure[17][5] , \gpio_configure[17][4] ,
         \gpio_configure[17][3] , \gpio_configure[17][2] ,
         \gpio_configure[17][1] , \gpio_configure[17][0] ,
         \gpio_configure[16][12] , \gpio_configure[16][11] ,
         \gpio_configure[16][10] , \gpio_configure[16][9] ,
         \gpio_configure[16][8] , \gpio_configure[16][7] ,
         \gpio_configure[16][6] , \gpio_configure[16][5] ,
         \gpio_configure[16][4] , \gpio_configure[16][3] ,
         \gpio_configure[16][2] , \gpio_configure[16][1] ,
         \gpio_configure[16][0] , \gpio_configure[15][12] ,
         \gpio_configure[15][11] , \gpio_configure[15][10] ,
         \gpio_configure[15][9] , \gpio_configure[15][8] ,
         \gpio_configure[15][7] , \gpio_configure[15][6] ,
         \gpio_configure[15][5] , \gpio_configure[15][4] ,
         \gpio_configure[15][3] , \gpio_configure[15][2] ,
         \gpio_configure[15][1] , \gpio_configure[15][0] ,
         \gpio_configure[14][12] , \gpio_configure[14][11] ,
         \gpio_configure[14][10] , \gpio_configure[14][9] ,
         \gpio_configure[14][8] , \gpio_configure[14][7] ,
         \gpio_configure[14][6] , \gpio_configure[14][5] ,
         \gpio_configure[14][4] , \gpio_configure[14][3] ,
         \gpio_configure[14][2] , \gpio_configure[14][1] ,
         \gpio_configure[14][0] , \gpio_configure[13][12] ,
         \gpio_configure[13][11] , \gpio_configure[13][10] ,
         \gpio_configure[13][9] , \gpio_configure[13][8] ,
         \gpio_configure[13][7] , \gpio_configure[13][6] ,
         \gpio_configure[13][5] , \gpio_configure[13][4] ,
         \gpio_configure[13][3] , \gpio_configure[13][2] ,
         \gpio_configure[13][1] , \gpio_configure[13][0] ,
         \gpio_configure[12][12] , \gpio_configure[12][11] ,
         \gpio_configure[12][10] , \gpio_configure[12][9] ,
         \gpio_configure[12][8] , \gpio_configure[12][7] ,
         \gpio_configure[12][6] , \gpio_configure[12][5] ,
         \gpio_configure[12][4] , \gpio_configure[12][3] ,
         \gpio_configure[12][2] , \gpio_configure[12][1] ,
         \gpio_configure[12][0] , \gpio_configure[11][12] ,
         \gpio_configure[11][11] , \gpio_configure[11][10] ,
         \gpio_configure[11][9] , \gpio_configure[11][8] ,
         \gpio_configure[11][7] , \gpio_configure[11][6] ,
         \gpio_configure[11][5] , \gpio_configure[11][4] ,
         \gpio_configure[11][3] , \gpio_configure[11][2] ,
         \gpio_configure[11][1] , \gpio_configure[11][0] ,
         \gpio_configure[10][12] , \gpio_configure[10][11] ,
         \gpio_configure[10][10] , \gpio_configure[10][9] ,
         \gpio_configure[10][8] , \gpio_configure[10][7] ,
         \gpio_configure[10][6] , \gpio_configure[10][5] ,
         \gpio_configure[10][4] , \gpio_configure[10][3] ,
         \gpio_configure[10][2] , \gpio_configure[10][1] ,
         \gpio_configure[10][0] , \gpio_configure[9][12] ,
         \gpio_configure[9][11] , \gpio_configure[9][10] ,
         \gpio_configure[9][9] , \gpio_configure[9][8] ,
         \gpio_configure[9][7] , \gpio_configure[9][6] ,
         \gpio_configure[9][5] , \gpio_configure[9][4] ,
         \gpio_configure[9][3] , \gpio_configure[9][2] ,
         \gpio_configure[9][1] , \gpio_configure[9][0] ,
         \gpio_configure[8][12] , \gpio_configure[8][11] ,
         \gpio_configure[8][10] , \gpio_configure[8][9] ,
         \gpio_configure[8][8] , \gpio_configure[8][7] ,
         \gpio_configure[8][6] , \gpio_configure[8][5] ,
         \gpio_configure[8][4] , \gpio_configure[8][3] ,
         \gpio_configure[8][2] , \gpio_configure[8][1] ,
         \gpio_configure[8][0] , \gpio_configure[7][12] ,
         \gpio_configure[7][11] , \gpio_configure[7][10] ,
         \gpio_configure[7][9] , \gpio_configure[7][8] ,
         \gpio_configure[7][7] , \gpio_configure[7][6] ,
         \gpio_configure[7][5] , \gpio_configure[7][4] ,
         \gpio_configure[7][3] , \gpio_configure[7][2] ,
         \gpio_configure[7][1] , \gpio_configure[7][0] ,
         \gpio_configure[6][12] , \gpio_configure[6][11] ,
         \gpio_configure[6][10] , \gpio_configure[6][9] ,
         \gpio_configure[6][8] , \gpio_configure[6][7] ,
         \gpio_configure[6][6] , \gpio_configure[6][5] ,
         \gpio_configure[6][4] , \gpio_configure[6][3] ,
         \gpio_configure[6][2] , \gpio_configure[6][1] ,
         \gpio_configure[6][0] , \gpio_configure[5][12] ,
         \gpio_configure[5][11] , \gpio_configure[5][10] ,
         \gpio_configure[5][9] , \gpio_configure[5][8] ,
         \gpio_configure[5][7] , \gpio_configure[5][6] ,
         \gpio_configure[5][5] , \gpio_configure[5][4] ,
         \gpio_configure[5][3] , \gpio_configure[5][2] ,
         \gpio_configure[5][1] , \gpio_configure[5][0] ,
         \gpio_configure[4][12] , \gpio_configure[4][11] ,
         \gpio_configure[4][10] , \gpio_configure[4][9] ,
         \gpio_configure[4][8] , \gpio_configure[4][7] ,
         \gpio_configure[4][6] , \gpio_configure[4][5] ,
         \gpio_configure[4][4] , \gpio_configure[4][3] ,
         \gpio_configure[4][2] , \gpio_configure[4][1] ,
         \gpio_configure[4][0] , \gpio_configure[3][12] ,
         \gpio_configure[3][11] , \gpio_configure[3][10] ,
         \gpio_configure[3][9] , \gpio_configure[3][8] ,
         \gpio_configure[3][7] , \gpio_configure[3][6] ,
         \gpio_configure[3][5] , \gpio_configure[3][4] ,
         \gpio_configure[3][3] , \gpio_configure[3][2] ,
         \gpio_configure[3][1] , \gpio_configure[3][0] ,
         \gpio_configure[2][12] , \gpio_configure[2][11] ,
         \gpio_configure[2][10] , \gpio_configure[2][9] ,
         \gpio_configure[2][8] , \gpio_configure[2][7] ,
         \gpio_configure[2][6] , \gpio_configure[2][5] ,
         \gpio_configure[2][4] , \gpio_configure[2][3] ,
         \gpio_configure[2][2] , \gpio_configure[2][1] ,
         \gpio_configure[2][0] , \gpio_configure[1][12] ,
         \gpio_configure[1][11] , \gpio_configure[1][10] ,
         \gpio_configure[1][9] , \gpio_configure[1][8] ,
         \gpio_configure[1][7] , \gpio_configure[1][6] ,
         \gpio_configure[1][5] , \gpio_configure[1][4] ,
         \gpio_configure[1][3] , \gpio_configure[1][2] ,
         \gpio_configure[1][1] , \gpio_configure[1][0] ,
         \gpio_configure[0][12] , \gpio_configure[0][11] ,
         \gpio_configure[0][10] , \gpio_configure[0][9] ,
         \gpio_configure[0][8] , \gpio_configure[0][7] ,
         \gpio_configure[0][6] , \gpio_configure[0][5] ,
         \gpio_configure[0][4] , \gpio_configure[0][3] ,
         \gpio_configure[0][2] , \gpio_configure[0][1] ,
         \gpio_configure[0][0] , hkspi_disable, spi_is_enabled, rdstb, wrstb,
         wbbd_sck, wbbd_write, wbbd_busy, N860, N861, N862, N863, N864, N865,
         N866, N867, N868, N869, \_1_net_[0] , sdo, sdo_enb, pass_thru_user,
         pass_thru_user_delay, mgmt_gpio_data_33, mgmt_gpio_data_32,
         mgmt_gpio_data_15, mgmt_gpio_data_14, mgmt_gpio_data_13,
         mgmt_gpio_data_10, mgmt_gpio_data_9, mgmt_gpio_data_8,
         mgmt_gpio_data_6, mgmt_gpio_data_1, mgmt_gpio_data_0,
         mgmt_gpio_out_9_prebuff, clk2_output_dest, mgmt_gpio_out_15_prebuff,
         clk1_output_dest, mgmt_gpio_out_14_prebuff, trap_output_dest,
         irq_1_inputsrc, irq_2_inputsrc, serial_bb_enable, serial_bb_clock,
         serial_clock_pre, serial_bb_resetn, serial_resetn_pre, serial_bb_load,
         serial_load_pre, serial_bb_data_1, serial_bb_data_2, serial_xfer,
         serial_busy, csclk, \hkspi/fixed[2] , \hkspi/fixed[1] ,
         \hkspi/fixed[0] , \hkspi/N34 , \hkspi/writemode , \hkspi/readmode ,
         \hkspi/count[2] , \hkspi/count[1] , \hkspi/count[0] ,
         \hkspi/pre_pass_thru_user , \hkspi/pre_pass_thru_mgmt ,
         \hkspi/ldata[6] , \hkspi/ldata[5] , \hkspi/ldata[4] ,
         \hkspi/ldata[3] , \hkspi/ldata[2] , \hkspi/ldata[1] ,
         \hkspi/ldata[0] , \hkspi/state[2] , \hkspi/state[1] ,
         \hkspi/state[0] , \hkspi/addr[7] , \hkspi/addr[6] , \hkspi/addr[5] ,
         \hkspi/addr[4] , \hkspi/addr[3] , \hkspi/addr[2] , \hkspi/addr[1] ,
         \hkspi/addr[0] , n386, n620, n633, n2319, n2322, n2335, n2340, n2341,
         n2342, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2320, n2321, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2336, n2337, n2338, n2339, n2343, n2535, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388;
  wire   [3:0] wbbd_state;
  wire   [7:0] wbbd_addr;
  wire   [7:0] wbbd_data;
  wire   [7:0] idata;
  wire   [37:35] mgmt_gpio_data;
  wire   [12:0] serial_data_staging_1;
  wire   [12:0] serial_data_staging_2;
  wire   [1:0] xfer_state;
  wire   [4:0] pad_count_1;
  wire   [5:0] pad_count_2;
  wire   [3:0] xfer_count;
  wire   [23:0] mgmt_gpio_data_buf;
  assign wb_rstn_i = wb_rstn_i_BAR;
  assign N860 = wb_adr_i[2];
  assign N861 = wb_adr_i[3];
  assign N862 = wb_adr_i[4];
  assign N863 = wb_adr_i[5];
  assign N864 = wb_adr_i[6];
  assign N865 = wb_adr_i[7];
  assign N866 = wb_adr_i[20];
  assign N867 = wb_adr_i[21];
  assign N868 = wb_adr_i[22];
  assign N869 = wb_adr_i[23];
  assign idata[0] = mgmt_gpio_in[2];
  assign mgmt_gpio_out[37] = mgmt_gpio_data[37];
  assign mgmt_gpio_out[36] = mgmt_gpio_data[36];
  assign mgmt_gpio_out[9] = mgmt_gpio_out_9_prebuff;
  assign mgmt_gpio_out[15] = mgmt_gpio_out_15_prebuff;
  assign mgmt_gpio_out[14] = mgmt_gpio_out_14_prebuff;

  dfcrq1 serial_resetn_pre_reg ( .D(1'b1), .CP(n3334), .CDN(n3387), .Q(
        serial_resetn_pre) );
  dfcrq1 \hkspi/fixed_reg[2]  ( .D(n3093), .CP(mgmt_gpio_in[4]), .CDN(n3295), 
        .Q(\hkspi/fixed[2] ) );
  dfcrq1 \hkspi/state_reg[1]  ( .D(n3096), .CP(n3291), .CDN(n3294), .Q(
        \hkspi/state[1] ) );
  dfcrq1 \hkspi/count_reg[1]  ( .D(n3098), .CP(n3291), .CDN(n3295), .Q(
        \hkspi/count[1] ) );
  dfcrq1 \hkspi/pre_pass_thru_mgmt_reg  ( .D(n3097), .CP(n3291), .CDN(n3295), 
        .Q(\hkspi/pre_pass_thru_mgmt ) );
  dfcrq1 \hkspi/state_reg[0]  ( .D(n3101), .CP(n3291), .CDN(n3294), .Q(
        \hkspi/state[0] ) );
  dfcrq1 \hkspi/pre_pass_thru_user_reg  ( .D(n3102), .CP(n3291), .CDN(n3294), 
        .Q(\hkspi/pre_pass_thru_user ) );
  dfcrq1 \hkspi/state_reg[2]  ( .D(n3103), .CP(n3291), .CDN(n3294), .Q(
        \hkspi/state[2] ) );
  dfcrq1 \hkspi/pass_thru_user_reg  ( .D(n3092), .CP(mgmt_gpio_in[4]), .CDN(
        n3294), .Q(pass_thru_user) );
  dfcrq1 \hkspi/pass_thru_mgmt_reg  ( .D(n3091), .CP(mgmt_gpio_in[4]), .CDN(
        n3294), .Q(pass_thru_mgmt) );
  dfcrq1 \hkspi/count_reg[0]  ( .D(n3100), .CP(mgmt_gpio_in[4]), .CDN(n3293), 
        .Q(\hkspi/count[0] ) );
  dfcrq1 \hkspi/count_reg[2]  ( .D(n3099), .CP(mgmt_gpio_in[4]), .CDN(n3294), 
        .Q(\hkspi/count[2] ) );
  dfcrq1 \hkspi/fixed_reg[0]  ( .D(n3095), .CP(mgmt_gpio_in[4]), .CDN(n3294), 
        .Q(\hkspi/fixed[0] ) );
  dfcrq1 \hkspi/fixed_reg[1]  ( .D(n3094), .CP(mgmt_gpio_in[4]), .CDN(n3294), 
        .Q(\hkspi/fixed[1] ) );
  dfcrq1 \hkspi/addr_reg[0]  ( .D(n3089), .CP(n3291), .CDN(n3294), .Q(
        \hkspi/addr[0] ) );
  dfcrq1 \hkspi/addr_reg[1]  ( .D(n3090), .CP(n3291), .CDN(n3293), .Q(
        \hkspi/addr[1] ) );
  dfcrq1 \hkspi/addr_reg[2]  ( .D(n3088), .CP(mgmt_gpio_in[4]), .CDN(n3293), 
        .Q(\hkspi/addr[2] ) );
  dfcrq1 \hkspi/addr_reg[3]  ( .D(n3087), .CP(mgmt_gpio_in[4]), .CDN(n3293), 
        .Q(\hkspi/addr[3] ) );
  dfcrq1 \hkspi/addr_reg[4]  ( .D(n3086), .CP(mgmt_gpio_in[4]), .CDN(n3293), 
        .Q(\hkspi/addr[4] ) );
  dfcrq1 \hkspi/addr_reg[5]  ( .D(n3085), .CP(mgmt_gpio_in[4]), .CDN(n3293), 
        .Q(\hkspi/addr[5] ) );
  dfcrq1 \hkspi/addr_reg[6]  ( .D(n3084), .CP(mgmt_gpio_in[4]), .CDN(n3293), 
        .Q(\hkspi/addr[6] ) );
  dfcrq1 \hkspi/addr_reg[7]  ( .D(n3083), .CP(mgmt_gpio_in[4]), .CDN(n3293), 
        .Q(\hkspi/addr[7] ) );
  dfcrq1 \hkspi/rdstb_reg  ( .D(n3082), .CP(mgmt_gpio_in[4]), .CDN(n3293), .Q(
        rdstb) );
  dfcrq1 \gpio_configure_reg[3][3]  ( .D(n2688), .CP(n3319), .CDN(n3383), .Q(
        \gpio_configure[3][3] ) );
  dfcrq1 \wbbd_state_reg[0]  ( .D(n3076), .CP(n3332), .CDN(n3388), .Q(
        wbbd_state[0]) );
  dfcrq1 \wbbd_state_reg[2]  ( .D(n3077), .CP(n3332), .CDN(n3388), .Q(
        wbbd_state[2]) );
  dfcrq1 \wbbd_state_reg[3]  ( .D(n3079), .CP(n3332), .CDN(n3388), .Q(
        wbbd_state[3]) );
  dfcrq1 \wbbd_state_reg[1]  ( .D(n3078), .CP(n3331), .CDN(n3388), .Q(
        wbbd_state[1]) );
  dfcrq1 \wbbd_addr_reg[0]  ( .D(n3067), .CP(n3331), .CDN(n3388), .Q(
        wbbd_addr[0]) );
  dfcrq1 \wbbd_addr_reg[1]  ( .D(n3066), .CP(n3331), .CDN(n3292), .Q(
        wbbd_addr[1]) );
  dfcrq1 \wbbd_addr_reg[2]  ( .D(n3065), .CP(n3331), .CDN(n3292), .Q(
        wbbd_addr[2]) );
  dfcrq1 \wbbd_addr_reg[3]  ( .D(n3064), .CP(n3331), .CDN(n3292), .Q(
        wbbd_addr[3]) );
  dfcrq1 \wbbd_addr_reg[4]  ( .D(n3063), .CP(n3331), .CDN(n3292), .Q(
        wbbd_addr[4]) );
  dfcrq1 \wbbd_addr_reg[5]  ( .D(n3062), .CP(n3331), .CDN(n3292), .Q(
        wbbd_addr[5]) );
  dfcrq1 \wbbd_addr_reg[6]  ( .D(n3061), .CP(n3331), .CDN(n3292), .Q(
        wbbd_addr[6]) );
  dfcrq1 \wbbd_data_reg[0]  ( .D(n3075), .CP(n3331), .CDN(n3292), .Q(
        wbbd_data[0]) );
  dfcrq1 \wbbd_data_reg[1]  ( .D(n3074), .CP(n3331), .CDN(n3292), .Q(
        wbbd_data[1]) );
  dfcrq1 \wbbd_data_reg[2]  ( .D(n3073), .CP(n3331), .CDN(n3292), .Q(
        wbbd_data[2]) );
  dfcrq1 \wbbd_data_reg[3]  ( .D(n3072), .CP(n3331), .CDN(n3292), .Q(
        wbbd_data[3]) );
  dfcrq1 \wbbd_data_reg[4]  ( .D(n3071), .CP(n3331), .CDN(n3292), .Q(
        wbbd_data[4]) );
  dfcrq1 \wbbd_data_reg[5]  ( .D(n3070), .CP(n3331), .CDN(n3292), .Q(
        wbbd_data[5]) );
  dfcrq1 \wbbd_data_reg[6]  ( .D(n3069), .CP(n3331), .CDN(n3292), .Q(
        wbbd_data[6]) );
  dfcrq1 \wbbd_data_reg[7]  ( .D(n3068), .CP(n3331), .CDN(n3292), .Q(
        wbbd_data[7]) );
  dfcrq1 wbbd_write_reg ( .D(n3059), .CP(n3334), .CDN(n3292), .Q(wbbd_write)
         );
  dfcrq1 wbbd_sck_reg ( .D(n3058), .CP(wb_clk_i), .CDN(n3292), .Q(wbbd_sck) );
  dfcrq1 \gpio_configure_reg[3][7]  ( .D(n2692), .CP(n3319), .CDN(n3375), .Q(
        \gpio_configure[3][7] ) );
  dfcrq1 \gpio_configure_reg[3][6]  ( .D(n2691), .CP(n3319), .CDN(n3387), .Q(
        \gpio_configure[3][6] ) );
  dfcrq1 \gpio_configure_reg[3][5]  ( .D(n2690), .CP(n3319), .CDN(n3383), .Q(
        \gpio_configure[3][5] ) );
  dfcrq1 \gpio_configure_reg[3][4]  ( .D(n2689), .CP(n3319), .CDN(n3375), .Q(
        \gpio_configure[3][4] ) );
  dfcrq1 \gpio_configure_reg[4][12]  ( .D(n2706), .CP(n3319), .CDN(porb), .Q(
        \gpio_configure[4][12] ) );
  dfcrq1 \gpio_configure_reg[4][11]  ( .D(n2705), .CP(n3319), .CDN(porb), .Q(
        \gpio_configure[4][11] ) );
  dfcrq1 \gpio_configure_reg[4][9]  ( .D(n2704), .CP(n3304), .CDN(porb), .Q(
        \gpio_configure[4][9] ) );
  dfcrq1 \gpio_configure_reg[4][8]  ( .D(n2703), .CP(n3304), .CDN(porb), .Q(
        \gpio_configure[4][8] ) );
  dfcrq1 \gpio_configure_reg[16][12]  ( .D(n2826), .CP(n3317), .CDN(porb), .Q(
        \gpio_configure[16][12] ) );
  dfcrq1 \gpio_configure_reg[16][11]  ( .D(n2825), .CP(n3322), .CDN(porb), .Q(
        \gpio_configure[16][11] ) );
  dfcrq1 \gpio_configure_reg[16][9]  ( .D(n2824), .CP(n3304), .CDN(n3386), .Q(
        \gpio_configure[16][9] ) );
  dfcrq1 \gpio_configure_reg[16][8]  ( .D(n2823), .CP(n3312), .CDN(n3382), .Q(
        \gpio_configure[16][8] ) );
  dfcrq1 \gpio_configure_reg[15][7]  ( .D(n2812), .CP(n3304), .CDN(n3381), .Q(
        \gpio_configure[15][7] ) );
  dfcrq1 \gpio_configure_reg[15][6]  ( .D(n2811), .CP(n3304), .CDN(n3386), .Q(
        \gpio_configure[15][6] ) );
  dfcrq1 \gpio_configure_reg[15][5]  ( .D(n2810), .CP(n3329), .CDN(n3382), .Q(
        \gpio_configure[15][5] ) );
  dfcrq1 \gpio_configure_reg[15][4]  ( .D(n2809), .CP(n3314), .CDN(n3381), .Q(
        \gpio_configure[15][4] ) );
  dfcrq1 \gpio_configure_reg[15][3]  ( .D(n2808), .CP(n3299), .CDN(n3386), .Q(
        \gpio_configure[15][3] ) );
  dfcrq1 \gpio_configure_reg[15][2]  ( .D(n2807), .CP(n3298), .CDN(n3382), .Q(
        \gpio_configure[15][2] ) );
  dfcrq1 \gpio_configure_reg[0][10]  ( .D(n2666), .CP(n3325), .CDN(n3381), .Q(
        \gpio_configure[0][10] ) );
  dfcrq1 \gpio_configure_reg[0][9]  ( .D(n2665), .CP(n3306), .CDN(n3386), .Q(
        \gpio_configure[0][9] ) );
  dfcrq1 \gpio_configure_reg[0][8]  ( .D(n2664), .CP(n3305), .CDN(n3385), .Q(
        \gpio_configure[0][8] ) );
  dfcrq1 irq_2_inputsrc_reg ( .D(n3056), .CP(n3329), .CDN(n3384), .Q(
        irq_2_inputsrc) );
  dfcrq1 irq_1_inputsrc_reg ( .D(n2601), .CP(n3302), .CDN(n3376), .Q(
        irq_1_inputsrc) );
  dfcrq1 \gpio_configure_reg[8][12]  ( .D(n2746), .CP(n3317), .CDN(n3385), .Q(
        \gpio_configure[8][12] ) );
  dfcrq1 \gpio_configure_reg[8][11]  ( .D(n2745), .CP(n3306), .CDN(n3384), .Q(
        \gpio_configure[8][11] ) );
  dfcrq1 \gpio_configure_reg[8][9]  ( .D(n2744), .CP(n3320), .CDN(n3376), .Q(
        \gpio_configure[8][9] ) );
  dfcrq1 \gpio_configure_reg[8][8]  ( .D(n2743), .CP(n3325), .CDN(n3385), .Q(
        \gpio_configure[8][8] ) );
  dfcrq1 \gpio_configure_reg[7][7]  ( .D(n2732), .CP(n3329), .CDN(n3384), .Q(
        \gpio_configure[7][7] ) );
  dfcrq1 \gpio_configure_reg[7][6]  ( .D(n2731), .CP(n3319), .CDN(n3376), .Q(
        \gpio_configure[7][6] ) );
  dfcrq1 \gpio_configure_reg[7][5]  ( .D(n2730), .CP(n3314), .CDN(n3385), .Q(
        \gpio_configure[7][5] ) );
  dfcrq1 \gpio_configure_reg[7][4]  ( .D(n2729), .CP(n3329), .CDN(n3384), .Q(
        \gpio_configure[7][4] ) );
  dfcrq1 \gpio_configure_reg[7][3]  ( .D(n2728), .CP(n3329), .CDN(n3376), .Q(
        \gpio_configure[7][3] ) );
  dfcrq1 \gpio_configure_reg[7][2]  ( .D(n2727), .CP(n3319), .CDN(n3385), .Q(
        \gpio_configure[7][2] ) );
  dfcrq1 \gpio_configure_reg[12][12]  ( .D(n2786), .CP(n3329), .CDN(n3384), 
        .Q(\gpio_configure[12][12] ) );
  dfcrq1 \gpio_configure_reg[12][11]  ( .D(n2785), .CP(n3314), .CDN(n3376), 
        .Q(\gpio_configure[12][11] ) );
  dfcrq1 \gpio_configure_reg[12][9]  ( .D(n2784), .CP(n3299), .CDN(n3385), .Q(
        \gpio_configure[12][9] ) );
  dfcrq1 \gpio_configure_reg[12][8]  ( .D(n2783), .CP(n3298), .CDN(n3384), .Q(
        \gpio_configure[12][8] ) );
  dfcrq1 \gpio_configure_reg[11][7]  ( .D(n2772), .CP(n3329), .CDN(n3376), .Q(
        \gpio_configure[11][7] ) );
  dfcrq1 \gpio_configure_reg[11][6]  ( .D(n2771), .CP(n3329), .CDN(n3385), .Q(
        \gpio_configure[11][6] ) );
  dfcrq1 \gpio_configure_reg[11][5]  ( .D(n2770), .CP(n3305), .CDN(n3384), .Q(
        \gpio_configure[11][5] ) );
  dfcrq1 \gpio_configure_reg[11][4]  ( .D(n2769), .CP(n3329), .CDN(n3375), .Q(
        \gpio_configure[11][4] ) );
  dfcrq1 \gpio_configure_reg[11][3]  ( .D(n2768), .CP(n3328), .CDN(n3387), .Q(
        \gpio_configure[11][3] ) );
  dfcrq1 \gpio_configure_reg[11][2]  ( .D(n2767), .CP(n3329), .CDN(n3383), .Q(
        \gpio_configure[11][2] ) );
  dfcrq1 \gpio_configure_reg[36][10]  ( .D(n3025), .CP(n3329), .CDN(n3375), 
        .Q(\gpio_configure[36][10] ) );
  dfcrq1 \gpio_configure_reg[36][9]  ( .D(n3024), .CP(n3319), .CDN(n3387), .Q(
        \gpio_configure[36][9] ) );
  dfcrq1 \gpio_configure_reg[36][8]  ( .D(n3023), .CP(n3319), .CDN(n3383), .Q(
        \gpio_configure[36][8] ) );
  dfcrq1 \gpio_configure_reg[35][7]  ( .D(n3012), .CP(n3318), .CDN(n3375), .Q(
        \gpio_configure[35][7] ) );
  dfcrq1 \gpio_configure_reg[35][6]  ( .D(n3011), .CP(n3318), .CDN(n3387), .Q(
        \gpio_configure[35][6] ) );
  dfcrq1 \gpio_configure_reg[35][5]  ( .D(n3010), .CP(n3318), .CDN(n3383), .Q(
        \gpio_configure[35][5] ) );
  dfcrq1 \gpio_configure_reg[35][4]  ( .D(n3009), .CP(n3318), .CDN(n3375), .Q(
        \gpio_configure[35][4] ) );
  dfcrq1 \gpio_configure_reg[35][3]  ( .D(n3008), .CP(n3318), .CDN(n3382), .Q(
        \gpio_configure[35][3] ) );
  dfcrq1 \gpio_configure_reg[35][2]  ( .D(n3007), .CP(n3318), .CDN(n3381), .Q(
        \gpio_configure[35][2] ) );
  dfcrq1 \gpio_configure_reg[20][12]  ( .D(n2866), .CP(n3318), .CDN(n3386), 
        .Q(\gpio_configure[20][12] ) );
  dfcrq1 \gpio_configure_reg[20][11]  ( .D(n2865), .CP(n3318), .CDN(n3382), 
        .Q(\gpio_configure[20][11] ) );
  dfcrq1 \gpio_configure_reg[20][9]  ( .D(n2864), .CP(n3328), .CDN(n3381), .Q(
        \gpio_configure[20][9] ) );
  dfcrq1 \gpio_configure_reg[20][8]  ( .D(n2863), .CP(n3318), .CDN(n3386), .Q(
        \gpio_configure[20][8] ) );
  dfcrq1 \gpio_configure_reg[19][7]  ( .D(n2852), .CP(n3308), .CDN(n3382), .Q(
        \gpio_configure[19][7] ) );
  dfcrq1 \gpio_configure_reg[19][6]  ( .D(n2851), .CP(n3328), .CDN(n3381), .Q(
        \gpio_configure[19][6] ) );
  dfcrq1 \gpio_configure_reg[19][5]  ( .D(n2850), .CP(n3318), .CDN(n3386), .Q(
        \gpio_configure[19][5] ) );
  dfcrq1 \gpio_configure_reg[19][4]  ( .D(n2849), .CP(n3327), .CDN(n3382), .Q(
        \gpio_configure[19][4] ) );
  dfcrq1 \gpio_configure_reg[19][3]  ( .D(n2848), .CP(n3323), .CDN(n3381), .Q(
        \gpio_configure[19][3] ) );
  dfcrq1 \gpio_configure_reg[19][2]  ( .D(n2847), .CP(n3328), .CDN(n3386), .Q(
        \gpio_configure[19][2] ) );
  dfcrq1 \gpio_configure_reg[24][12]  ( .D(n2906), .CP(n3318), .CDN(n3382), 
        .Q(\gpio_configure[24][12] ) );
  dfcrq1 \gpio_configure_reg[24][11]  ( .D(n2905), .CP(n3318), .CDN(n3381), 
        .Q(\gpio_configure[24][11] ) );
  dfcrq1 \gpio_configure_reg[24][9]  ( .D(n2904), .CP(n3328), .CDN(n3386), .Q(
        \gpio_configure[24][9] ) );
  dfcrq1 \gpio_configure_reg[24][8]  ( .D(n2903), .CP(n3318), .CDN(n3382), .Q(
        \gpio_configure[24][8] ) );
  dfcrq1 \gpio_configure_reg[23][7]  ( .D(n2892), .CP(n3327), .CDN(n3381), .Q(
        \gpio_configure[23][7] ) );
  dfcrq1 \gpio_configure_reg[23][6]  ( .D(n2891), .CP(n3328), .CDN(n3386), .Q(
        \gpio_configure[23][6] ) );
  dfcrq1 \gpio_configure_reg[23][5]  ( .D(n2890), .CP(n3307), .CDN(n3382), .Q(
        \gpio_configure[23][5] ) );
  dfcrq1 \gpio_configure_reg[23][4]  ( .D(n2889), .CP(n3318), .CDN(n3381), .Q(
        \gpio_configure[23][4] ) );
  dfcrq1 \gpio_configure_reg[23][3]  ( .D(n2888), .CP(n3313), .CDN(n3380), .Q(
        \gpio_configure[23][3] ) );
  dfcrq1 \gpio_configure_reg[23][2]  ( .D(n2887), .CP(n3319), .CDN(n3380), .Q(
        \gpio_configure[23][2] ) );
  dfcrq1 \gpio_configure_reg[32][12]  ( .D(n2986), .CP(n3312), .CDN(n3380), 
        .Q(\gpio_configure[32][12] ) );
  dfcrq1 \gpio_configure_reg[32][11]  ( .D(n2985), .CP(n3317), .CDN(n3380), 
        .Q(\gpio_configure[32][11] ) );
  dfcrq1 \gpio_configure_reg[32][9]  ( .D(n2984), .CP(n3315), .CDN(n3380), .Q(
        \gpio_configure[32][9] ) );
  dfcrq1 \gpio_configure_reg[32][8]  ( .D(n2983), .CP(n3312), .CDN(n3380), .Q(
        \gpio_configure[32][8] ) );
  dfcrq1 \gpio_configure_reg[31][7]  ( .D(n2972), .CP(n3313), .CDN(n3380), .Q(
        \gpio_configure[31][7] ) );
  dfcrq1 \gpio_configure_reg[31][6]  ( .D(n2971), .CP(n3320), .CDN(n3380), .Q(
        \gpio_configure[31][6] ) );
  dfcrq1 \gpio_configure_reg[31][5]  ( .D(n2970), .CP(n3328), .CDN(n3380), .Q(
        \gpio_configure[31][5] ) );
  dfcrq1 \gpio_configure_reg[31][4]  ( .D(n2969), .CP(n3328), .CDN(n3380), .Q(
        \gpio_configure[31][4] ) );
  dfcrq1 \gpio_configure_reg[31][3]  ( .D(n2968), .CP(n3328), .CDN(n3337), .Q(
        \gpio_configure[31][3] ) );
  dfcrq1 \gpio_configure_reg[31][2]  ( .D(n2967), .CP(n3318), .CDN(n3336), .Q(
        \gpio_configure[31][2] ) );
  dfcrq1 \gpio_configure_reg[28][12]  ( .D(n2946), .CP(n3328), .CDN(n3338), 
        .Q(\gpio_configure[28][12] ) );
  dfcrq1 \gpio_configure_reg[28][11]  ( .D(n2945), .CP(n3328), .CDN(n3339), 
        .Q(\gpio_configure[28][11] ) );
  dfcrq1 \gpio_configure_reg[28][9]  ( .D(n2944), .CP(n3328), .CDN(n3337), .Q(
        \gpio_configure[28][9] ) );
  dfcrq1 \gpio_configure_reg[28][8]  ( .D(n2943), .CP(n3327), .CDN(n3336), .Q(
        \gpio_configure[28][8] ) );
  dfcrq1 \gpio_configure_reg[27][7]  ( .D(n2932), .CP(n3328), .CDN(n3338), .Q(
        \gpio_configure[27][7] ) );
  dfcrq1 \gpio_configure_reg[27][6]  ( .D(n2931), .CP(n3328), .CDN(n3339), .Q(
        \gpio_configure[27][6] ) );
  dfcrq1 \gpio_configure_reg[27][5]  ( .D(n2930), .CP(n3328), .CDN(n3337), .Q(
        \gpio_configure[27][5] ) );
  dfcrq1 \gpio_configure_reg[27][4]  ( .D(n2929), .CP(n3318), .CDN(n3336), .Q(
        \gpio_configure[27][4] ) );
  dfcrq1 \gpio_configure_reg[27][3]  ( .D(n2928), .CP(n3328), .CDN(n3378), .Q(
        \gpio_configure[27][3] ) );
  dfcrq1 \gpio_configure_reg[27][2]  ( .D(n2927), .CP(n3328), .CDN(n3378), .Q(
        \gpio_configure[27][2] ) );
  dfcrq1 serial_xfer_reg ( .D(n3055), .CP(n3323), .CDN(n3378), .Q(serial_xfer)
         );
  dfcrq1 serial_bb_enable_reg ( .D(n3040), .CP(n3323), .CDN(n3378), .Q(
        serial_bb_enable) );
  dfcrq1 serial_bb_data_2_reg ( .D(n3039), .CP(n3308), .CDN(n3378), .Q(
        serial_bb_data_2) );
  dfcrq1 serial_bb_data_1_reg ( .D(n3038), .CP(n3307), .CDN(n3378), .Q(
        serial_bb_data_1) );
  dfcrq1 serial_bb_clock_reg ( .D(n3037), .CP(n3305), .CDN(n3378), .Q(
        serial_bb_clock) );
  dfcrq1 \xfer_count_reg[0]  ( .D(n2628), .CP(n3333), .CDN(n3378), .Q(
        xfer_count[0]) );
  dfcrq1 \xfer_count_reg[2]  ( .D(n2626), .CP(n3332), .CDN(n3378), .Q(
        xfer_count[2]) );
  dfcrq1 \xfer_state_reg[1]  ( .D(n2655), .CP(n3331), .CDN(n3387), .Q(
        xfer_state[1]) );
  dfcrq1 \xfer_state_reg[0]  ( .D(n2656), .CP(n3330), .CDN(n3377), .Q(
        xfer_state[0]) );
  dfcrq1 \xfer_count_reg[1]  ( .D(n2627), .CP(n3334), .CDN(n3377), .Q(
        xfer_count[1]) );
  dfcrq1 \xfer_count_reg[3]  ( .D(n2629), .CP(n3334), .CDN(n3377), .Q(
        xfer_count[3]) );
  dfcrq1 serial_load_pre_reg ( .D(n2624), .CP(n3334), .CDN(n3377), .Q(
        serial_load_pre) );
  dfcrq1 \pad_count_2_reg[2]  ( .D(n2622), .CP(wb_clk_i), .CDN(n3377), .Q(
        pad_count_2[2]) );
  dfcrq1 \pad_count_2_reg[3]  ( .D(n2621), .CP(n3334), .CDN(n3377), .Q(
        pad_count_2[3]) );
  dfcrq1 \pad_count_2_reg[5]  ( .D(n2620), .CP(wb_clk_i), .CDN(n3377), .Q(
        pad_count_2[5]) );
  dfcrq1 \pad_count_1_reg[0]  ( .D(n2619), .CP(wb_clk_i), .CDN(n3377), .Q(
        pad_count_1[0]) );
  dfcrq1 \pad_count_1_reg[2]  ( .D(n2618), .CP(n3334), .CDN(n3377), .Q(
        pad_count_1[2]) );
  dfcrq1 \pad_count_1_reg[3]  ( .D(n2617), .CP(n3330), .CDN(n3377), .Q(
        pad_count_1[3]) );
  dfcrq1 serial_busy_reg ( .D(n2623), .CP(n3330), .CDN(n3376), .Q(serial_busy)
         );
  dfcrq1 serial_clock_pre_reg ( .D(n2625), .CP(n3330), .CDN(n3385), .Q(
        serial_clock_pre) );
  dfcrq1 serial_bb_load_reg ( .D(n3036), .CP(n3308), .CDN(n3384), .Q(
        serial_bb_load) );
  dfcrq1 serial_bb_resetn_reg ( .D(n3035), .CP(n3307), .CDN(n3376), .Q(
        serial_bb_resetn) );
  dfcrq1 \gpio_configure_reg[11][12]  ( .D(n2776), .CP(n3305), .CDN(n3385), 
        .Q(\gpio_configure[11][12] ) );
  dfcrq1 \gpio_configure_reg[11][11]  ( .D(n2775), .CP(n3327), .CDN(n3384), 
        .Q(\gpio_configure[11][11] ) );
  dfcrq1 \gpio_configure_reg[11][9]  ( .D(n2774), .CP(n3308), .CDN(n3376), .Q(
        \gpio_configure[11][9] ) );
  dfcrq1 \gpio_configure_reg[11][8]  ( .D(n2773), .CP(n3308), .CDN(n3385), .Q(
        \gpio_configure[11][8] ) );
  dfcrq1 \gpio_configure_reg[10][7]  ( .D(n2762), .CP(n3307), .CDN(n3384), .Q(
        \gpio_configure[10][7] ) );
  dfcrq1 \gpio_configure_reg[10][6]  ( .D(n2761), .CP(n3305), .CDN(n3376), .Q(
        \gpio_configure[10][6] ) );
  dfcrq1 \gpio_configure_reg[10][5]  ( .D(n2760), .CP(n3306), .CDN(n3383), .Q(
        \gpio_configure[10][5] ) );
  dfcrq1 \gpio_configure_reg[10][4]  ( .D(n2759), .CP(n3327), .CDN(n3375), .Q(
        \gpio_configure[10][4] ) );
  dfcrq1 \gpio_configure_reg[10][3]  ( .D(n2758), .CP(n3305), .CDN(n3387), .Q(
        \gpio_configure[10][3] ) );
  dfcrq1 \gpio_configure_reg[10][2]  ( .D(n2757), .CP(n3308), .CDN(n3383), .Q(
        \gpio_configure[10][2] ) );
  dfcrq1 \pll_div_reg[4]  ( .D(n2611), .CP(n3307), .CDN(n3375), .Q(pll_div[4])
         );
  dfcrq1 \pll_div_reg[3]  ( .D(n2610), .CP(n3305), .CDN(n3387), .Q(pll_div[3])
         );
  dfcrq1 \pll_div_reg[1]  ( .D(n2609), .CP(n3306), .CDN(n3383), .Q(pll_div[1])
         );
  dfcrq1 \pll_div_reg[0]  ( .D(n2608), .CP(n3327), .CDN(n3375), .Q(pll_div[0])
         );
  dfcrq1 \gpio_configure_reg[3][12]  ( .D(n2696), .CP(n3323), .CDN(n3387), .Q(
        \gpio_configure[3][12] ) );
  dfcrq1 \gpio_configure_reg[3][10]  ( .D(n2695), .CP(n3327), .CDN(n3383), .Q(
        \gpio_configure[3][10] ) );
  dfcrq1 \gpio_configure_reg[3][9]  ( .D(n2694), .CP(n3323), .CDN(n3368), .Q(
        \gpio_configure[3][9] ) );
  dfcrq1 \gpio_configure_reg[3][8]  ( .D(n2693), .CP(n3323), .CDN(n3372), .Q(
        \gpio_configure[3][8] ) );
  dfcrq1 \gpio_configure_reg[7][12]  ( .D(n2736), .CP(n3307), .CDN(n3368), .Q(
        \gpio_configure[7][12] ) );
  dfcrq1 \gpio_configure_reg[7][11]  ( .D(n2735), .CP(n3310), .CDN(n3369), .Q(
        \gpio_configure[7][11] ) );
  dfcrq1 \gpio_configure_reg[7][9]  ( .D(n2734), .CP(n3323), .CDN(n3369), .Q(
        \gpio_configure[7][9] ) );
  dfcrq1 \gpio_configure_reg[7][8]  ( .D(n2733), .CP(csclk), .CDN(n3371), .Q(
        \gpio_configure[7][8] ) );
  dfcrq1 \gpio_configure_reg[6][7]  ( .D(n2722), .CP(csclk), .CDN(n3368), .Q(
        \gpio_configure[6][7] ) );
  dfcrq1 \gpio_configure_reg[6][6]  ( .D(n2721), .CP(csclk), .CDN(n3369), .Q(
        \gpio_configure[6][6] ) );
  dfcrq1 \gpio_configure_reg[6][5]  ( .D(n2720), .CP(n3309), .CDN(n3371), .Q(
        \gpio_configure[6][5] ) );
  dfcrq1 \gpio_configure_reg[6][4]  ( .D(n2719), .CP(n3310), .CDN(n3369), .Q(
        \gpio_configure[6][4] ) );
  dfcrq1 \gpio_configure_reg[6][3]  ( .D(n2718), .CP(n3304), .CDN(n3374), .Q(
        \gpio_configure[6][3] ) );
  dfcrq1 \gpio_configure_reg[6][2]  ( .D(n2717), .CP(n3327), .CDN(n3370), .Q(
        \gpio_configure[6][2] ) );
  dfcrq1 irq_spi_reg ( .D(n2606), .CP(n3327), .CDN(n3368), .Q(irq[0]) );
  dfcrq1 reset_reg_reg ( .D(n2605), .CP(n3323), .CDN(n3369), .Q(reset_reg) );
  dfcrq1 \gpio_configure_reg[15][12]  ( .D(n2816), .CP(n3305), .CDN(n3370), 
        .Q(\gpio_configure[15][12] ) );
  dfcrq1 \gpio_configure_reg[15][11]  ( .D(n2815), .CP(n3308), .CDN(n3368), 
        .Q(\gpio_configure[15][11] ) );
  dfcrq1 \gpio_configure_reg[15][9]  ( .D(n2814), .CP(n3307), .CDN(n3372), .Q(
        \gpio_configure[15][9] ) );
  dfcrq1 \gpio_configure_reg[15][8]  ( .D(n2813), .CP(n3305), .CDN(n3373), .Q(
        \gpio_configure[15][8] ) );
  dfcrq1 \gpio_configure_reg[14][7]  ( .D(n2802), .CP(n3306), .CDN(n3374), .Q(
        \gpio_configure[14][7] ) );
  dfcrq1 \gpio_configure_reg[14][6]  ( .D(n2801), .CP(n3327), .CDN(n3369), .Q(
        \gpio_configure[14][6] ) );
  dfcrq1 \gpio_configure_reg[14][5]  ( .D(n2800), .CP(n3327), .CDN(n3370), .Q(
        \gpio_configure[14][5] ) );
  dfcrq1 \gpio_configure_reg[14][4]  ( .D(n2799), .CP(n3327), .CDN(n3371), .Q(
        \gpio_configure[14][4] ) );
  dfcrq1 \gpio_configure_reg[14][3]  ( .D(n2798), .CP(n3327), .CDN(n3374), .Q(
        \gpio_configure[14][3] ) );
  dfcrq1 \gpio_configure_reg[14][2]  ( .D(n2797), .CP(n3327), .CDN(n3370), .Q(
        \gpio_configure[14][2] ) );
  dfcrq1 clk1_output_dest_reg ( .D(n2604), .CP(n3308), .CDN(n3372), .Q(
        clk1_output_dest) );
  dfcrq1 clk2_output_dest_reg ( .D(n2603), .CP(n3308), .CDN(n3373), .Q(
        clk2_output_dest) );
  dfcrq1 trap_output_dest_reg ( .D(n2602), .CP(n3307), .CDN(n3370), .Q(
        trap_output_dest) );
  dfcrq1 \gpio_configure_reg[35][12]  ( .D(n3016), .CP(n3317), .CDN(n3371), 
        .Q(\gpio_configure[35][12] ) );
  dfcrq1 \gpio_configure_reg[35][11]  ( .D(n3015), .CP(n3317), .CDN(n3368), 
        .Q(\gpio_configure[35][11] ) );
  dfcrq1 \gpio_configure_reg[35][9]  ( .D(n3014), .CP(n3317), .CDN(n3370), .Q(
        \gpio_configure[35][9] ) );
  dfcrq1 \gpio_configure_reg[35][8]  ( .D(n3013), .CP(n3317), .CDN(n3368), .Q(
        \gpio_configure[35][8] ) );
  dfcrq1 \gpio_configure_reg[34][7]  ( .D(n3002), .CP(n3317), .CDN(n3373), .Q(
        \gpio_configure[34][7] ) );
  dfcrq1 \gpio_configure_reg[34][6]  ( .D(n3001), .CP(n3317), .CDN(n3370), .Q(
        \gpio_configure[34][6] ) );
  dfcrq1 \gpio_configure_reg[34][5]  ( .D(n3000), .CP(n3317), .CDN(n3371), .Q(
        \gpio_configure[34][5] ) );
  dfcrq1 \gpio_configure_reg[34][4]  ( .D(n2999), .CP(n3317), .CDN(n3373), .Q(
        \gpio_configure[34][4] ) );
  dfcrq1 \gpio_configure_reg[34][3]  ( .D(n2998), .CP(n3316), .CDN(n3371), .Q(
        \gpio_configure[34][3] ) );
  dfcrq1 \gpio_configure_reg[34][2]  ( .D(n2997), .CP(n3316), .CDN(n3370), .Q(
        \gpio_configure[34][2] ) );
  dfcrq1 \gpio_configure_reg[19][12]  ( .D(n2856), .CP(n3316), .CDN(n3371), 
        .Q(\gpio_configure[19][12] ) );
  dfcrq1 \gpio_configure_reg[19][11]  ( .D(n2855), .CP(n3316), .CDN(n3372), 
        .Q(\gpio_configure[19][11] ) );
  dfcrq1 \gpio_configure_reg[19][9]  ( .D(n2854), .CP(n3316), .CDN(n3371), .Q(
        \gpio_configure[19][9] ) );
  dfcrq1 \gpio_configure_reg[19][8]  ( .D(n2853), .CP(n3316), .CDN(n3374), .Q(
        \gpio_configure[19][8] ) );
  dfcrq1 \gpio_configure_reg[18][7]  ( .D(n2842), .CP(n3316), .CDN(n3371), .Q(
        \gpio_configure[18][7] ) );
  dfcrq1 \gpio_configure_reg[18][6]  ( .D(n2841), .CP(n3316), .CDN(n3372), .Q(
        \gpio_configure[18][6] ) );
  dfcrq1 \gpio_configure_reg[18][5]  ( .D(n2840), .CP(n3315), .CDN(n3374), .Q(
        \gpio_configure[18][5] ) );
  dfcrq1 \gpio_configure_reg[18][4]  ( .D(n2839), .CP(n3315), .CDN(n3368), .Q(
        \gpio_configure[18][4] ) );
  dfcrq1 \gpio_configure_reg[18][3]  ( .D(n2838), .CP(n3315), .CDN(n3370), .Q(
        \gpio_configure[18][3] ) );
  dfcrq1 \gpio_configure_reg[18][2]  ( .D(n2837), .CP(n3315), .CDN(n3369), .Q(
        \gpio_configure[18][2] ) );
  dfcrq1 \gpio_configure_reg[23][12]  ( .D(n2896), .CP(n3315), .CDN(n3373), 
        .Q(\gpio_configure[23][12] ) );
  dfcrq1 \gpio_configure_reg[23][11]  ( .D(n2895), .CP(n3315), .CDN(n3368), 
        .Q(\gpio_configure[23][11] ) );
  dfcrq1 \gpio_configure_reg[23][9]  ( .D(n2894), .CP(n3315), .CDN(n3371), .Q(
        \gpio_configure[23][9] ) );
  dfcrq1 \gpio_configure_reg[23][8]  ( .D(n2893), .CP(n3315), .CDN(n3373), .Q(
        \gpio_configure[23][8] ) );
  dfcrq1 \gpio_configure_reg[22][7]  ( .D(n2882), .CP(n3314), .CDN(n3369), .Q(
        \gpio_configure[22][7] ) );
  dfcrq1 \gpio_configure_reg[22][6]  ( .D(n2881), .CP(n3314), .CDN(n3369), .Q(
        \gpio_configure[22][6] ) );
  dfcrq1 \gpio_configure_reg[22][5]  ( .D(n2880), .CP(n3314), .CDN(n3370), .Q(
        \gpio_configure[22][5] ) );
  dfcrq1 \gpio_configure_reg[22][4]  ( .D(n2879), .CP(n3314), .CDN(n3372), .Q(
        \gpio_configure[22][4] ) );
  dfcrq1 \gpio_configure_reg[22][3]  ( .D(n2878), .CP(n3314), .CDN(n3369), .Q(
        \gpio_configure[22][3] ) );
  dfcrq1 \gpio_configure_reg[22][2]  ( .D(n2877), .CP(n3314), .CDN(n3368), .Q(
        \gpio_configure[22][2] ) );
  dfcrq1 \gpio_configure_reg[31][12]  ( .D(n2976), .CP(n3314), .CDN(n3372), 
        .Q(\gpio_configure[31][12] ) );
  dfcrq1 \gpio_configure_reg[31][11]  ( .D(n2975), .CP(n3314), .CDN(n3368), 
        .Q(\gpio_configure[31][11] ) );
  dfcrq1 \gpio_configure_reg[31][9]  ( .D(n2974), .CP(n3313), .CDN(n3370), .Q(
        \gpio_configure[31][9] ) );
  dfcrq1 \gpio_configure_reg[31][8]  ( .D(n2973), .CP(n3313), .CDN(n3374), .Q(
        \gpio_configure[31][8] ) );
  dfcrq1 \gpio_configure_reg[30][7]  ( .D(n2962), .CP(n3313), .CDN(n3371), .Q(
        \gpio_configure[30][7] ) );
  dfcrq1 \gpio_configure_reg[30][6]  ( .D(n2961), .CP(n3313), .CDN(n3370), .Q(
        \gpio_configure[30][6] ) );
  dfcrq1 \gpio_configure_reg[30][5]  ( .D(n2960), .CP(n3313), .CDN(n3369), .Q(
        \gpio_configure[30][5] ) );
  dfcrq1 \gpio_configure_reg[30][4]  ( .D(n2959), .CP(n3313), .CDN(n3370), .Q(
        \gpio_configure[30][4] ) );
  dfcrq1 \gpio_configure_reg[30][3]  ( .D(n2958), .CP(n3313), .CDN(n3369), .Q(
        \gpio_configure[30][3] ) );
  dfcrq1 \gpio_configure_reg[30][2]  ( .D(n2957), .CP(n3313), .CDN(n3371), .Q(
        \gpio_configure[30][2] ) );
  dfcrq1 \gpio_configure_reg[27][12]  ( .D(n2936), .CP(n3312), .CDN(n3373), 
        .Q(\gpio_configure[27][12] ) );
  dfcrq1 \gpio_configure_reg[27][11]  ( .D(n2935), .CP(n3312), .CDN(n3368), 
        .Q(\gpio_configure[27][11] ) );
  dfcrq1 \gpio_configure_reg[27][9]  ( .D(n2934), .CP(n3312), .CDN(n3374), .Q(
        \gpio_configure[27][9] ) );
  dfcrq1 \gpio_configure_reg[27][8]  ( .D(n2933), .CP(n3312), .CDN(n3366), .Q(
        \gpio_configure[27][8] ) );
  dfcrq1 \gpio_configure_reg[26][7]  ( .D(n2922), .CP(n3312), .CDN(n3363), .Q(
        \gpio_configure[26][7] ) );
  dfcrq1 \gpio_configure_reg[26][6]  ( .D(n2921), .CP(n3312), .CDN(n3362), .Q(
        \gpio_configure[26][6] ) );
  dfcrq1 \gpio_configure_reg[26][5]  ( .D(n2920), .CP(n3312), .CDN(n3366), .Q(
        \gpio_configure[26][5] ) );
  dfcrq1 \gpio_configure_reg[26][4]  ( .D(n2919), .CP(n3312), .CDN(n3367), .Q(
        \gpio_configure[26][4] ) );
  dfcrq1 \gpio_configure_reg[26][3]  ( .D(n2918), .CP(n3311), .CDN(n3361), .Q(
        \gpio_configure[26][3] ) );
  dfcrq1 \gpio_configure_reg[26][2]  ( .D(n2917), .CP(n3311), .CDN(n3366), .Q(
        \gpio_configure[26][2] ) );
  dfcrq1 \gpio_configure_reg[14][12]  ( .D(n2806), .CP(n3311), .CDN(n3363), 
        .Q(\gpio_configure[14][12] ) );
  dfcrq1 \gpio_configure_reg[14][11]  ( .D(n2805), .CP(n3311), .CDN(n3364), 
        .Q(\gpio_configure[14][11] ) );
  dfcrq1 \gpio_configure_reg[14][9]  ( .D(n2804), .CP(n3311), .CDN(n3366), .Q(
        \gpio_configure[14][9] ) );
  dfcrq1 \gpio_configure_reg[14][8]  ( .D(n2803), .CP(n3311), .CDN(n3362), .Q(
        \gpio_configure[14][8] ) );
  dfcrq1 \gpio_configure_reg[13][7]  ( .D(n2792), .CP(n3311), .CDN(n3363), .Q(
        \gpio_configure[13][7] ) );
  dfcrq1 \gpio_configure_reg[13][6]  ( .D(n2791), .CP(n3311), .CDN(n3367), .Q(
        \gpio_configure[13][6] ) );
  dfcrq1 \gpio_configure_reg[13][5]  ( .D(n2790), .CP(n3311), .CDN(n3362), .Q(
        \gpio_configure[13][5] ) );
  dfcrq1 \gpio_configure_reg[13][4]  ( .D(n2789), .CP(n3305), .CDN(n3364), .Q(
        \gpio_configure[13][4] ) );
  dfcrq1 \gpio_configure_reg[13][3]  ( .D(n2788), .CP(n3327), .CDN(n3366), .Q(
        \gpio_configure[13][3] ) );
  dfcrq1 \gpio_configure_reg[13][2]  ( .D(n2787), .CP(n3326), .CDN(n3365), .Q(
        \gpio_configure[13][2] ) );
  dfcrq1 \gpio_configure_reg[10][12]  ( .D(n2766), .CP(n3311), .CDN(n3361), 
        .Q(\gpio_configure[10][12] ) );
  dfcrq1 \gpio_configure_reg[10][11]  ( .D(n2765), .CP(n3327), .CDN(n3364), 
        .Q(\gpio_configure[10][11] ) );
  dfcrq1 \gpio_configure_reg[10][9]  ( .D(n2764), .CP(n3326), .CDN(n3363), .Q(
        \gpio_configure[10][9] ) );
  dfcrq1 \gpio_configure_reg[10][8]  ( .D(n2763), .CP(n3311), .CDN(n3361), .Q(
        \gpio_configure[10][8] ) );
  dfcrq1 \gpio_configure_reg[9][7]  ( .D(n2752), .CP(n3311), .CDN(n3365), .Q(
        \gpio_configure[9][7] ) );
  dfcrq1 \gpio_configure_reg[9][6]  ( .D(n2751), .CP(n3326), .CDN(n3365), .Q(
        \gpio_configure[9][6] ) );
  dfcrq1 \gpio_configure_reg[9][5]  ( .D(n2750), .CP(n3326), .CDN(n3366), .Q(
        \gpio_configure[9][5] ) );
  dfcrq1 \gpio_configure_reg[9][4]  ( .D(n2749), .CP(n3311), .CDN(n3367), .Q(
        \gpio_configure[9][4] ) );
  dfcrq1 \gpio_configure_reg[9][3]  ( .D(n2748), .CP(n3311), .CDN(n3365), .Q(
        \gpio_configure[9][3] ) );
  dfcrq1 \gpio_configure_reg[9][2]  ( .D(n2747), .CP(n3326), .CDN(n3364), .Q(
        \gpio_configure[9][2] ) );
  dfcrq1 \pll_sel_reg[2]  ( .D(n2615), .CP(n3311), .CDN(n3367), .Q(pll_sel[2])
         );
  dfcrq1 \pll_sel_reg[0]  ( .D(n2614), .CP(n3326), .CDN(n3364), .Q(pll_sel[0])
         );
  dfcrq1 \pll90_sel_reg[2]  ( .D(n2613), .CP(n3325), .CDN(n3366), .Q(
        pll90_sel[2]) );
  dfcrq1 \pll90_sel_reg[0]  ( .D(n2612), .CP(n3329), .CDN(n3362), .Q(
        pll90_sel[0]) );
  dfcrq1 \gpio_configure_reg[6][12]  ( .D(n2726), .CP(n3319), .CDN(n3363), .Q(
        \gpio_configure[6][12] ) );
  dfcrq1 \gpio_configure_reg[6][11]  ( .D(n2725), .CP(n3314), .CDN(n3366), .Q(
        \gpio_configure[6][11] ) );
  dfcrq1 \gpio_configure_reg[6][9]  ( .D(n2724), .CP(n3312), .CDN(n3365), .Q(
        \gpio_configure[6][9] ) );
  dfcrq1 \gpio_configure_reg[6][8]  ( .D(n2723), .CP(n3309), .CDN(n3366), .Q(
        \gpio_configure[6][8] ) );
  dfcrq1 \gpio_configure_reg[5][7]  ( .D(n2712), .CP(n3317), .CDN(n3365), .Q(
        \gpio_configure[5][7] ) );
  dfcrq1 \gpio_configure_reg[5][6]  ( .D(n2711), .CP(n3318), .CDN(n3363), .Q(
        \gpio_configure[5][6] ) );
  dfcrq1 \gpio_configure_reg[5][5]  ( .D(n2710), .CP(n3326), .CDN(n3361), .Q(
        \gpio_configure[5][5] ) );
  dfcrq1 \gpio_configure_reg[5][4]  ( .D(n2709), .CP(n3326), .CDN(n3364), .Q(
        \gpio_configure[5][4] ) );
  dfcrq1 \gpio_configure_reg[5][3]  ( .D(n2708), .CP(n3326), .CDN(n3362), .Q(
        \gpio_configure[5][3] ) );
  dfcrq1 \gpio_configure_reg[5][2]  ( .D(n2707), .CP(n3311), .CDN(n3364), .Q(
        \gpio_configure[5][2] ) );
  dfcrq1 pll_ena_reg ( .D(n2607), .CP(n3326), .CDN(n3361), .Q(pll_ena) );
  dfcrq1 \gpio_configure_reg[2][12]  ( .D(n2685), .CP(n3326), .CDN(n3366), .Q(
        \gpio_configure[2][12] ) );
  dfcrq1 \gpio_configure_reg[2][11]  ( .D(n2684), .CP(n3326), .CDN(n3363), .Q(
        \gpio_configure[2][11] ) );
  dfcrq1 \gpio_configure_reg[2][9]  ( .D(n2683), .CP(n3326), .CDN(n3361), .Q(
        \gpio_configure[2][9] ) );
  dfcrq1 \gpio_configure_reg[2][8]  ( .D(n2682), .CP(n3326), .CDN(n3363), .Q(
        \gpio_configure[2][8] ) );
  dfcrq1 \mgmt_gpio_data_reg[37]  ( .D(n3054), .CP(n3326), .CDN(n3366), .Q(
        mgmt_gpio_data[37]) );
  dfcrq1 \mgmt_gpio_data_reg[36]  ( .D(n3053), .CP(n3311), .CDN(n3363), .Q(
        mgmt_gpio_data[36]) );
  dfcrq1 \mgmt_gpio_data_reg[35]  ( .D(n3052), .CP(n3326), .CDN(n3367), .Q(
        mgmt_gpio_data[35]) );
  dfcrq1 \mgmt_gpio_data_reg[34]  ( .D(n3051), .CP(n3326), .CDN(n3363), .Q(
        mgmt_gpio_out[34]) );
  dfcrq1 \mgmt_gpio_data_reg[33]  ( .D(n3050), .CP(n3326), .CDN(n3364), .Q(
        mgmt_gpio_data_33) );
  dfcrq1 \mgmt_gpio_data_reg[32]  ( .D(n3049), .CP(n3311), .CDN(n3367), .Q(
        mgmt_gpio_data_32) );
  dfcrq1 \gpio_configure_reg[37][7]  ( .D(n3031), .CP(n3311), .CDN(n3364), .Q(
        \gpio_configure[37][7] ) );
  dfcrq1 \gpio_configure_reg[37][6]  ( .D(n3030), .CP(n3310), .CDN(n3365), .Q(
        \gpio_configure[37][6] ) );
  dfcrq1 \gpio_configure_reg[37][5]  ( .D(n3029), .CP(n3310), .CDN(n3365), .Q(
        \gpio_configure[37][5] ) );
  dfcrq1 \gpio_configure_reg[37][4]  ( .D(n3028), .CP(n3310), .CDN(n3363), .Q(
        \gpio_configure[37][4] ) );
  dfcrq1 \gpio_configure_reg[37][3]  ( .D(n3027), .CP(n3310), .CDN(n3364), .Q(
        \gpio_configure[37][3] ) );
  dfcrq1 \gpio_configure_reg[37][2]  ( .D(n3026), .CP(n3310), .CDN(n3365), .Q(
        \gpio_configure[37][2] ) );
  dfcrq1 \gpio_configure_reg[22][12]  ( .D(n2886), .CP(n3310), .CDN(n3363), 
        .Q(\gpio_configure[22][12] ) );
  dfcrq1 \gpio_configure_reg[22][11]  ( .D(n2885), .CP(n3310), .CDN(n3365), 
        .Q(\gpio_configure[22][11] ) );
  dfcrq1 \gpio_configure_reg[22][9]  ( .D(n2884), .CP(n3310), .CDN(n3362), .Q(
        \gpio_configure[22][9] ) );
  dfcrq1 \gpio_configure_reg[22][8]  ( .D(n2883), .CP(n3309), .CDN(n3366), .Q(
        \gpio_configure[22][8] ) );
  dfcrq1 \gpio_configure_reg[21][7]  ( .D(n2872), .CP(n3309), .CDN(n3364), .Q(
        \gpio_configure[21][7] ) );
  dfcrq1 \gpio_configure_reg[21][6]  ( .D(n2871), .CP(n3309), .CDN(n3365), .Q(
        \gpio_configure[21][6] ) );
  dfcrq1 \gpio_configure_reg[21][5]  ( .D(n2870), .CP(n3309), .CDN(n3366), .Q(
        \gpio_configure[21][5] ) );
  dfcrq1 \gpio_configure_reg[21][4]  ( .D(n2869), .CP(n3309), .CDN(n3364), .Q(
        \gpio_configure[21][4] ) );
  dfcrq1 \gpio_configure_reg[21][3]  ( .D(n2868), .CP(n3309), .CDN(n3367), .Q(
        \gpio_configure[21][3] ) );
  dfcrq1 \gpio_configure_reg[21][2]  ( .D(n2867), .CP(n3309), .CDN(n3361), .Q(
        \gpio_configure[21][2] ) );
  dfcrq1 \gpio_configure_reg[34][12]  ( .D(n3006), .CP(n3309), .CDN(n3362), 
        .Q(\gpio_configure[34][12] ) );
  dfcrq1 \gpio_configure_reg[34][11]  ( .D(n3005), .CP(n3310), .CDN(n3365), 
        .Q(\gpio_configure[34][11] ) );
  dfcrq1 \gpio_configure_reg[34][9]  ( .D(n3004), .CP(n3309), .CDN(n3354), .Q(
        \gpio_configure[34][9] ) );
  dfcrq1 \gpio_configure_reg[34][8]  ( .D(n3003), .CP(n3325), .CDN(n3358), .Q(
        \gpio_configure[34][8] ) );
  dfcrq1 \gpio_configure_reg[33][7]  ( .D(n2992), .CP(n3310), .CDN(n3356), .Q(
        \gpio_configure[33][7] ) );
  dfcrq1 \gpio_configure_reg[33][6]  ( .D(n2991), .CP(n3309), .CDN(n3357), .Q(
        \gpio_configure[33][6] ) );
  dfcrq1 \gpio_configure_reg[33][5]  ( .D(n2990), .CP(n3325), .CDN(n3358), .Q(
        \gpio_configure[33][5] ) );
  dfcrq1 \gpio_configure_reg[33][4]  ( .D(n2989), .CP(n3310), .CDN(n3356), .Q(
        \gpio_configure[33][4] ) );
  dfcrq1 \gpio_configure_reg[33][3]  ( .D(n2988), .CP(n3309), .CDN(n3359), .Q(
        \gpio_configure[33][3] ) );
  dfcrq1 \gpio_configure_reg[33][2]  ( .D(n2987), .CP(n3319), .CDN(n3360), .Q(
        \gpio_configure[33][2] ) );
  dfcrq1 \gpio_configure_reg[18][12]  ( .D(n2846), .CP(csclk), .CDN(n3354), 
        .Q(\gpio_configure[18][12] ) );
  dfcrq1 \gpio_configure_reg[18][11]  ( .D(n2845), .CP(n3306), .CDN(n3357), 
        .Q(\gpio_configure[18][11] ) );
  dfcrq1 \gpio_configure_reg[18][9]  ( .D(n2844), .CP(n3316), .CDN(n3358), .Q(
        \gpio_configure[18][9] ) );
  dfcrq1 \gpio_configure_reg[18][8]  ( .D(n2843), .CP(n3320), .CDN(n3355), .Q(
        \gpio_configure[18][8] ) );
  dfcrq1 \gpio_configure_reg[17][7]  ( .D(n2832), .CP(csclk), .CDN(n3354), .Q(
        \gpio_configure[17][7] ) );
  dfcrq1 \gpio_configure_reg[17][6]  ( .D(n2831), .CP(n3329), .CDN(n3358), .Q(
        \gpio_configure[17][6] ) );
  dfcrq1 \gpio_configure_reg[17][5]  ( .D(n2830), .CP(n3319), .CDN(n3359), .Q(
        \gpio_configure[17][5] ) );
  dfcrq1 \gpio_configure_reg[17][4]  ( .D(n2829), .CP(n3325), .CDN(n3360), .Q(
        \gpio_configure[17][4] ) );
  dfcrq1 \gpio_configure_reg[17][3]  ( .D(n2828), .CP(n3325), .CDN(n3358), .Q(
        \gpio_configure[17][3] ) );
  dfcrq1 \gpio_configure_reg[17][2]  ( .D(n2827), .CP(n3325), .CDN(n3355), .Q(
        \gpio_configure[17][2] ) );
  dfcrq1 \gpio_configure_reg[30][12]  ( .D(n2966), .CP(n3310), .CDN(n3356), 
        .Q(\gpio_configure[30][12] ) );
  dfcrq1 \gpio_configure_reg[30][11]  ( .D(n2965), .CP(n3309), .CDN(n3358), 
        .Q(\gpio_configure[30][11] ) );
  dfcrq1 \gpio_configure_reg[30][9]  ( .D(n2964), .CP(n3325), .CDN(n3354), .Q(
        \gpio_configure[30][9] ) );
  dfcrq1 \gpio_configure_reg[30][8]  ( .D(n2963), .CP(n3325), .CDN(n3355), .Q(
        \gpio_configure[30][8] ) );
  dfcrq1 \gpio_configure_reg[29][7]  ( .D(n2952), .CP(n3325), .CDN(n3359), .Q(
        \gpio_configure[29][7] ) );
  dfcrq1 \gpio_configure_reg[29][6]  ( .D(n2951), .CP(n3325), .CDN(n3354), .Q(
        \gpio_configure[29][6] ) );
  dfcrq1 \gpio_configure_reg[29][5]  ( .D(n2950), .CP(n3325), .CDN(n3356), .Q(
        \gpio_configure[29][5] ) );
  dfcrq1 \gpio_configure_reg[29][4]  ( .D(n2949), .CP(n3310), .CDN(n3358), .Q(
        \gpio_configure[29][4] ) );
  dfcrq1 \gpio_configure_reg[29][3]  ( .D(n2948), .CP(n3309), .CDN(n3357), .Q(
        \gpio_configure[29][3] ) );
  dfcrq1 \gpio_configure_reg[29][2]  ( .D(n2947), .CP(n3325), .CDN(n3360), .Q(
        \gpio_configure[29][2] ) );
  dfcrq1 \gpio_configure_reg[26][12]  ( .D(n2926), .CP(n3325), .CDN(n3356), 
        .Q(\gpio_configure[26][12] ) );
  dfcrq1 \gpio_configure_reg[26][11]  ( .D(n2925), .CP(n3310), .CDN(n3355), 
        .Q(\gpio_configure[26][11] ) );
  dfcrq1 \gpio_configure_reg[26][9]  ( .D(n2924), .CP(n3309), .CDN(n3360), .Q(
        \gpio_configure[26][9] ) );
  dfcrq1 \gpio_configure_reg[26][8]  ( .D(n2923), .CP(n3308), .CDN(n3357), .Q(
        \gpio_configure[26][8] ) );
  dfcrq1 \gpio_configure_reg[25][7]  ( .D(n2912), .CP(n3308), .CDN(n3357), .Q(
        \gpio_configure[25][7] ) );
  dfcrq1 \gpio_configure_reg[25][6]  ( .D(n2911), .CP(n3308), .CDN(n3358), .Q(
        \gpio_configure[25][6] ) );
  dfcrq1 \gpio_configure_reg[25][5]  ( .D(n2910), .CP(n3308), .CDN(n3359), .Q(
        \gpio_configure[25][5] ) );
  dfcrq1 \gpio_configure_reg[25][4]  ( .D(n2909), .CP(n3308), .CDN(n3357), .Q(
        \gpio_configure[25][4] ) );
  dfcrq1 \gpio_configure_reg[25][3]  ( .D(n2908), .CP(n3308), .CDN(n3356), .Q(
        \gpio_configure[25][3] ) );
  dfcrq1 \gpio_configure_reg[25][2]  ( .D(n2907), .CP(n3308), .CDN(n3359), .Q(
        \gpio_configure[25][2] ) );
  dfcrq1 \gpio_configure_reg[5][12]  ( .D(n2716), .CP(n3308), .CDN(n3356), .Q(
        \gpio_configure[5][12] ) );
  dfcrq1 \gpio_configure_reg[5][11]  ( .D(n2715), .CP(n3312), .CDN(n3358), .Q(
        \gpio_configure[5][11] ) );
  dfcrq1 \gpio_configure_reg[5][9]  ( .D(n2714), .CP(n3312), .CDN(n3354), .Q(
        \gpio_configure[5][9] ) );
  dfcrq1 \gpio_configure_reg[5][8]  ( .D(n2713), .CP(n3312), .CDN(n3355), .Q(
        \gpio_configure[5][8] ) );
  dfcrq1 \gpio_configure_reg[4][7]  ( .D(n2702), .CP(n3312), .CDN(n3358), .Q(
        \gpio_configure[4][7] ) );
  dfcrq1 \gpio_configure_reg[4][6]  ( .D(n2701), .CP(n3312), .CDN(n3357), .Q(
        \gpio_configure[4][6] ) );
  dfcrq1 \gpio_configure_reg[4][5]  ( .D(n2700), .CP(n3312), .CDN(n3358), .Q(
        \gpio_configure[4][5] ) );
  dfcrq1 \gpio_configure_reg[4][4]  ( .D(n2699), .CP(n3312), .CDN(n3357), .Q(
        \gpio_configure[4][4] ) );
  dfcrq1 \gpio_configure_reg[4][3]  ( .D(n2698), .CP(n3312), .CDN(n3355), .Q(
        \gpio_configure[4][3] ) );
  dfcrq1 \gpio_configure_reg[4][2]  ( .D(n2697), .CP(n3307), .CDN(n3360), .Q(
        \gpio_configure[4][2] ) );
  dfcrq1 \gpio_configure_reg[13][12]  ( .D(n2796), .CP(n3307), .CDN(n3356), 
        .Q(\gpio_configure[13][12] ) );
  dfcrq1 \gpio_configure_reg[13][11]  ( .D(n2795), .CP(n3307), .CDN(n3354), 
        .Q(\gpio_configure[13][11] ) );
  dfcrq1 \gpio_configure_reg[13][9]  ( .D(n2794), .CP(n3307), .CDN(n3356), .Q(
        \gpio_configure[13][9] ) );
  dfcrq1 \gpio_configure_reg[13][8]  ( .D(n2793), .CP(n3307), .CDN(n3360), .Q(
        \gpio_configure[13][8] ) );
  dfcrq1 \gpio_configure_reg[12][7]  ( .D(n2782), .CP(n3307), .CDN(n3358), .Q(
        \gpio_configure[12][7] ) );
  dfcrq1 \gpio_configure_reg[12][6]  ( .D(n2781), .CP(n3307), .CDN(n3355), .Q(
        \gpio_configure[12][6] ) );
  dfcrq1 \gpio_configure_reg[12][5]  ( .D(n2780), .CP(n3307), .CDN(n3360), .Q(
        \gpio_configure[12][5] ) );
  dfcrq1 \gpio_configure_reg[12][4]  ( .D(n2779), .CP(n3322), .CDN(n3355), .Q(
        \gpio_configure[12][4] ) );
  dfcrq1 \gpio_configure_reg[12][3]  ( .D(n2778), .CP(n3314), .CDN(n3358), .Q(
        \gpio_configure[12][3] ) );
  dfcrq1 \gpio_configure_reg[12][2]  ( .D(n2777), .CP(n3316), .CDN(n3355), .Q(
        \gpio_configure[12][2] ) );
  dfcrq1 \gpio_configure_reg[17][12]  ( .D(n2836), .CP(csclk), .CDN(n3359), 
        .Q(\gpio_configure[17][12] ) );
  dfcrq1 \gpio_configure_reg[17][11]  ( .D(n2835), .CP(n3303), .CDN(n3355), 
        .Q(\gpio_configure[17][11] ) );
  dfcrq1 \gpio_configure_reg[17][9]  ( .D(n2834), .CP(n3320), .CDN(n3356), .Q(
        \gpio_configure[17][9] ) );
  dfcrq1 \gpio_configure_reg[17][8]  ( .D(n2833), .CP(n3306), .CDN(n3359), .Q(
        \gpio_configure[17][8] ) );
  dfcrq1 \gpio_configure_reg[16][7]  ( .D(n2822), .CP(csclk), .CDN(n3356), .Q(
        \gpio_configure[16][7] ) );
  dfcrq1 \gpio_configure_reg[16][6]  ( .D(n2821), .CP(n3306), .CDN(n3357), .Q(
        \gpio_configure[16][6] ) );
  dfcrq1 \gpio_configure_reg[16][5]  ( .D(n2820), .CP(n3306), .CDN(n3357), .Q(
        \gpio_configure[16][5] ) );
  dfcrq1 \gpio_configure_reg[16][4]  ( .D(n2819), .CP(n3306), .CDN(n3355), .Q(
        \gpio_configure[16][4] ) );
  dfcrq1 \gpio_configure_reg[16][3]  ( .D(n2818), .CP(n3306), .CDN(n3356), .Q(
        \gpio_configure[16][3] ) );
  dfcrq1 \gpio_configure_reg[16][2]  ( .D(n2817), .CP(n3306), .CDN(n3357), .Q(
        \gpio_configure[16][2] ) );
  dfcrq1 \gpio_configure_reg[1][10]  ( .D(n2675), .CP(n3306), .CDN(n3355), .Q(
        \gpio_configure[1][10] ) );
  dfcrq1 \gpio_configure_reg[1][9]  ( .D(n2674), .CP(n3306), .CDN(n3357), .Q(
        \gpio_configure[1][9] ) );
  dfcrq1 \gpio_configure_reg[1][8]  ( .D(n2673), .CP(n3306), .CDN(n3349), .Q(
        \gpio_configure[1][8] ) );
  dfcrq1 \gpio_configure_reg[0][7]  ( .D(n2663), .CP(n3305), .CDN(n3352), .Q(
        \gpio_configure[0][7] ) );
  dfcrq1 \gpio_configure_reg[0][6]  ( .D(n2662), .CP(n3305), .CDN(n3349), .Q(
        \gpio_configure[0][6] ) );
  dfcrq1 \gpio_configure_reg[0][5]  ( .D(n2661), .CP(n3305), .CDN(n3350), .Q(
        \gpio_configure[0][5] ) );
  dfcrq1 \gpio_configure_reg[0][4]  ( .D(n2660), .CP(n3305), .CDN(n3350), .Q(
        \gpio_configure[0][4] ) );
  dfcrq1 \gpio_configure_reg[0][3]  ( .D(n2659), .CP(n3305), .CDN(n3348), .Q(
        \gpio_configure[0][3] ) );
  dfcrq1 \gpio_configure_reg[0][2]  ( .D(n2658), .CP(n3305), .CDN(n3349), .Q(
        \gpio_configure[0][2] ) );
  dfcrq1 \gpio_configure_reg[9][12]  ( .D(n2756), .CP(n3305), .CDN(n3350), .Q(
        \gpio_configure[9][12] ) );
  dfcrq1 \gpio_configure_reg[9][11]  ( .D(n2755), .CP(n3305), .CDN(n3348), .Q(
        \gpio_configure[9][11] ) );
  dfcrq1 \gpio_configure_reg[9][9]  ( .D(n2754), .CP(n3304), .CDN(n3350), .Q(
        \gpio_configure[9][9] ) );
  dfcrq1 \gpio_configure_reg[9][8]  ( .D(n2753), .CP(n3304), .CDN(porb), .Q(
        \gpio_configure[9][8] ) );
  dfcrq1 \gpio_configure_reg[8][7]  ( .D(n2742), .CP(n3304), .CDN(n3351), .Q(
        \gpio_configure[8][7] ) );
  dfcrq1 \gpio_configure_reg[8][6]  ( .D(n2741), .CP(n3304), .CDN(n3349), .Q(
        \gpio_configure[8][6] ) );
  dfcrq1 \gpio_configure_reg[8][5]  ( .D(n2740), .CP(n3304), .CDN(n3350), .Q(
        \gpio_configure[8][5] ) );
  dfcrq1 \gpio_configure_reg[8][4]  ( .D(n2739), .CP(n3304), .CDN(n3351), .Q(
        \gpio_configure[8][4] ) );
  dfcrq1 \gpio_configure_reg[8][3]  ( .D(n2738), .CP(n3304), .CDN(n3349), .Q(
        \gpio_configure[8][3] ) );
  dfcrq1 \gpio_configure_reg[8][2]  ( .D(n2737), .CP(n3304), .CDN(n3352), .Q(
        \gpio_configure[8][2] ) );
  dfcrq1 \pll_trim_reg[12]  ( .D(n2616), .CP(n3303), .CDN(n3353), .Q(
        pll_trim[12]) );
  dfcrq1 hkspi_disable_reg ( .D(n3080), .CP(n3303), .CDN(n3339), .Q(
        hkspi_disable) );
  dfcrq1 \gpio_configure_reg[25][12]  ( .D(n2916), .CP(n3303), .CDN(n3350), 
        .Q(\gpio_configure[25][12] ) );
  dfcrq1 \gpio_configure_reg[25][11]  ( .D(n2915), .CP(n3303), .CDN(n3351), 
        .Q(\gpio_configure[25][11] ) );
  dfcrq1 \gpio_configure_reg[25][9]  ( .D(n2914), .CP(n3303), .CDN(n3348), .Q(
        \gpio_configure[25][9] ) );
  dfcrq1 \gpio_configure_reg[25][8]  ( .D(n2913), .CP(n3303), .CDN(n3343), .Q(
        \gpio_configure[25][8] ) );
  dfcrq1 \gpio_configure_reg[24][7]  ( .D(n2902), .CP(n3303), .CDN(n3351), .Q(
        \gpio_configure[24][7] ) );
  dfcrq1 \gpio_configure_reg[24][6]  ( .D(n2901), .CP(n3303), .CDN(n3352), .Q(
        \gpio_configure[24][6] ) );
  dfcrq1 \gpio_configure_reg[24][5]  ( .D(n2900), .CP(n3302), .CDN(n3353), .Q(
        \gpio_configure[24][5] ) );
  dfcrq1 \gpio_configure_reg[24][4]  ( .D(n2899), .CP(n3302), .CDN(n3351), .Q(
        \gpio_configure[24][4] ) );
  dfcrq1 \gpio_configure_reg[24][3]  ( .D(n2898), .CP(n3302), .CDN(n3348), .Q(
        \gpio_configure[24][3] ) );
  dfcrq1 \gpio_configure_reg[24][2]  ( .D(n2897), .CP(n3302), .CDN(n3349), .Q(
        \gpio_configure[24][2] ) );
  dfcrq1 \gpio_configure_reg[37][10]  ( .D(n3034), .CP(n3302), .CDN(n3351), 
        .Q(\gpio_configure[37][10] ) );
  dfcrq1 \gpio_configure_reg[37][9]  ( .D(n3033), .CP(n3302), .CDN(porb), .Q(
        \gpio_configure[37][9] ) );
  dfcrq1 \gpio_configure_reg[37][8]  ( .D(n3032), .CP(n3302), .CDN(n3348), .Q(
        \gpio_configure[37][8] ) );
  dfcrq1 \gpio_configure_reg[36][7]  ( .D(n3022), .CP(n3302), .CDN(n3352), .Q(
        \gpio_configure[36][7] ) );
  dfcrq1 \gpio_configure_reg[36][6]  ( .D(n3021), .CP(n3314), .CDN(n3338), .Q(
        \gpio_configure[36][6] ) );
  dfcrq1 \gpio_configure_reg[36][5]  ( .D(n3020), .CP(n3299), .CDN(n3349), .Q(
        \gpio_configure[36][5] ) );
  dfcrq1 \gpio_configure_reg[36][4]  ( .D(n3019), .CP(n3298), .CDN(n3351), .Q(
        \gpio_configure[36][4] ) );
  dfcrq1 \gpio_configure_reg[36][3]  ( .D(n3018), .CP(n3306), .CDN(n3350), .Q(
        \gpio_configure[36][3] ) );
  dfcrq1 \gpio_configure_reg[36][2]  ( .D(n3017), .CP(n3314), .CDN(n3353), .Q(
        \gpio_configure[36][2] ) );
  dfcrq1 \gpio_configure_reg[21][12]  ( .D(n2876), .CP(n3321), .CDN(n3349), 
        .Q(\gpio_configure[21][12] ) );
  dfcrq1 \gpio_configure_reg[21][11]  ( .D(n2875), .CP(n3329), .CDN(n3348), 
        .Q(\gpio_configure[21][11] ) );
  dfcrq1 \gpio_configure_reg[21][9]  ( .D(n2874), .CP(n3319), .CDN(n3353), .Q(
        \gpio_configure[21][9] ) );
  dfcrq1 \gpio_configure_reg[21][8]  ( .D(n2873), .CP(n3304), .CDN(n3350), .Q(
        \gpio_configure[21][8] ) );
  dfcrq1 \gpio_configure_reg[20][7]  ( .D(n2862), .CP(n3298), .CDN(n3350), .Q(
        \gpio_configure[20][7] ) );
  dfcrq1 \gpio_configure_reg[20][6]  ( .D(n2861), .CP(n3317), .CDN(n3351), .Q(
        \gpio_configure[20][6] ) );
  dfcrq1 \gpio_configure_reg[20][5]  ( .D(n2860), .CP(n3313), .CDN(n3352), .Q(
        \gpio_configure[20][5] ) );
  dfcrq1 \gpio_configure_reg[20][4]  ( .D(n2859), .CP(n3299), .CDN(n3350), .Q(
        \gpio_configure[20][4] ) );
  dfcrq1 \gpio_configure_reg[20][3]  ( .D(n2858), .CP(n3315), .CDN(n3349), .Q(
        \gpio_configure[20][3] ) );
  dfcrq1 \gpio_configure_reg[20][2]  ( .D(n2857), .CP(n3302), .CDN(n3352), .Q(
        \gpio_configure[20][2] ) );
  dfcrq1 \gpio_configure_reg[33][12]  ( .D(n2996), .CP(n3316), .CDN(n3349), 
        .Q(\gpio_configure[33][12] ) );
  dfcrq1 \gpio_configure_reg[33][11]  ( .D(n2995), .CP(n3301), .CDN(n3351), 
        .Q(\gpio_configure[33][11] ) );
  dfcrq1 \gpio_configure_reg[33][9]  ( .D(n2994), .CP(n3301), .CDN(n3379), .Q(
        \gpio_configure[33][9] ) );
  dfcrq1 \gpio_configure_reg[33][8]  ( .D(n2993), .CP(n3301), .CDN(n3348), .Q(
        \gpio_configure[33][8] ) );
  dfcrq1 \gpio_configure_reg[32][7]  ( .D(n2982), .CP(n3301), .CDN(n3351), .Q(
        \gpio_configure[32][7] ) );
  dfcrq1 \gpio_configure_reg[32][6]  ( .D(n2981), .CP(n3301), .CDN(n3350), .Q(
        \gpio_configure[32][6] ) );
  dfcrq1 \gpio_configure_reg[32][5]  ( .D(n2980), .CP(n3301), .CDN(n3351), .Q(
        \gpio_configure[32][5] ) );
  dfcrq1 \gpio_configure_reg[32][4]  ( .D(n2979), .CP(n3301), .CDN(n3350), .Q(
        \gpio_configure[32][4] ) );
  dfcrq1 \gpio_configure_reg[32][3]  ( .D(n2978), .CP(n3301), .CDN(n3348), .Q(
        \gpio_configure[32][3] ) );
  dfcrq1 \gpio_configure_reg[32][2]  ( .D(n2977), .CP(n3300), .CDN(n3353), .Q(
        \gpio_configure[32][2] ) );
  dfcrq1 \gpio_configure_reg[29][12]  ( .D(n2956), .CP(n3300), .CDN(n3349), 
        .Q(\gpio_configure[29][12] ) );
  dfcrq1 \gpio_configure_reg[29][11]  ( .D(n2955), .CP(n3300), .CDN(porb), .Q(
        \gpio_configure[29][11] ) );
  dfcrq1 \gpio_configure_reg[29][9]  ( .D(n2954), .CP(n3300), .CDN(n3349), .Q(
        \gpio_configure[29][9] ) );
  dfcrq1 \gpio_configure_reg[29][8]  ( .D(n2953), .CP(n3300), .CDN(n3353), .Q(
        \gpio_configure[29][8] ) );
  dfcrq1 \gpio_configure_reg[28][7]  ( .D(n2942), .CP(n3300), .CDN(n3351), .Q(
        \gpio_configure[28][7] ) );
  dfcrq1 \gpio_configure_reg[28][6]  ( .D(n2941), .CP(n3300), .CDN(n3348), .Q(
        \gpio_configure[28][6] ) );
  dfcrq1 \gpio_configure_reg[28][5]  ( .D(n2940), .CP(n3300), .CDN(n3353), .Q(
        \gpio_configure[28][5] ) );
  dfcrq1 \gpio_configure_reg[28][4]  ( .D(n2939), .CP(n3324), .CDN(n3348), .Q(
        \gpio_configure[28][4] ) );
  dfcrq1 \gpio_configure_reg[28][3]  ( .D(n2938), .CP(n3300), .CDN(n3351), .Q(
        \gpio_configure[28][3] ) );
  dfcrq1 \gpio_configure_reg[28][2]  ( .D(n2937), .CP(n3321), .CDN(n3348), .Q(
        \gpio_configure[28][2] ) );
  dfcrq1 wb_ack_o_reg ( .D(n3057), .CP(n3330), .CDN(n3292), .Q(wb_ack_o) );
  dfcrq1 \gpio_configure_reg[3][2]  ( .D(n2687), .CP(n3321), .CDN(n3352), .Q(
        \gpio_configure[3][2] ) );
  dfcrq1 \gpio_configure_reg[3][1]  ( .D(n2686), .CP(n3324), .CDN(n3348), .Q(
        \gpio_configure[3][1] ) );
  dfcrq1 \gpio_configure_reg[2][7]  ( .D(n2681), .CP(n3300), .CDN(n3349), .Q(
        \gpio_configure[2][7] ) );
  dfcrq1 \gpio_configure_reg[2][6]  ( .D(n2680), .CP(n3321), .CDN(n3387), .Q(
        \gpio_configure[2][6] ) );
  dfcrq1 \gpio_configure_reg[2][5]  ( .D(n2679), .CP(n3324), .CDN(n3336), .Q(
        \gpio_configure[2][5] ) );
  dfcrq1 \gpio_configure_reg[2][4]  ( .D(n2678), .CP(n3321), .CDN(n3376), .Q(
        \gpio_configure[2][4] ) );
  dfcrq1 \gpio_configure_reg[2][3]  ( .D(n2677), .CP(n3300), .CDN(n3343), .Q(
        \gpio_configure[2][3] ) );
  dfcrq1 \gpio_configure_reg[2][2]  ( .D(n2676), .CP(n3324), .CDN(n3381), .Q(
        \gpio_configure[2][2] ) );
  dfcrq1 \gpio_configure_reg[1][7]  ( .D(n2672), .CP(n3324), .CDN(n3378), .Q(
        \gpio_configure[1][7] ) );
  dfcrq1 \gpio_configure_reg[1][6]  ( .D(n2671), .CP(n3300), .CDN(n3336), .Q(
        \gpio_configure[1][6] ) );
  dfcrq1 \gpio_configure_reg[1][5]  ( .D(n2670), .CP(n3300), .CDN(n3386), .Q(
        \gpio_configure[1][5] ) );
  dfcrq1 \gpio_configure_reg[1][4]  ( .D(n2669), .CP(n3324), .CDN(n3383), .Q(
        \gpio_configure[1][4] ) );
  dfcrq1 \gpio_configure_reg[1][3]  ( .D(n2668), .CP(n3300), .CDN(n3384), .Q(
        \gpio_configure[1][3] ) );
  dfcrq1 \gpio_configure_reg[1][2]  ( .D(n2667), .CP(n3302), .CDN(n3368), .Q(
        \gpio_configure[1][2] ) );
  dfcrq1 \serial_data_staging_1_reg[0]  ( .D(n2654), .CP(n3330), .CDN(n3343), 
        .Q(serial_data_staging_1[0]) );
  dfcrq1 \serial_data_staging_1_reg[1]  ( .D(n2653), .CP(n3330), .CDN(n3350), 
        .Q(serial_data_staging_1[1]) );
  dfcrq1 \serial_data_staging_1_reg[2]  ( .D(n2652), .CP(n3330), .CDN(n3356), 
        .Q(serial_data_staging_1[2]) );
  dfcrq1 \serial_data_staging_1_reg[3]  ( .D(n2651), .CP(n3330), .CDN(n3337), 
        .Q(serial_data_staging_1[3]) );
  dfcrq1 \serial_data_staging_1_reg[4]  ( .D(n2650), .CP(n3330), .CDN(n3339), 
        .Q(serial_data_staging_1[4]) );
  dfcrq1 \serial_data_staging_1_reg[5]  ( .D(n2649), .CP(n3330), .CDN(n3375), 
        .Q(serial_data_staging_1[5]) );
  dfcrq1 \serial_data_staging_1_reg[6]  ( .D(n2648), .CP(n3330), .CDN(n3378), 
        .Q(serial_data_staging_1[6]) );
  dfcrq1 \serial_data_staging_1_reg[7]  ( .D(n2647), .CP(n3330), .CDN(n3339), 
        .Q(serial_data_staging_1[7]) );
  dfcrq1 \serial_data_staging_1_reg[8]  ( .D(n2646), .CP(n3330), .CDN(n3364), 
        .Q(serial_data_staging_1[8]) );
  dfcrq1 \serial_data_staging_1_reg[9]  ( .D(n2645), .CP(n3330), .CDN(n3376), 
        .Q(serial_data_staging_1[9]) );
  dfcrq1 \serial_data_staging_1_reg[10]  ( .D(n2644), .CP(n3330), .CDN(n3387), 
        .Q(serial_data_staging_1[10]) );
  dfcrq1 \serial_data_staging_1_reg[11]  ( .D(n2643), .CP(n3330), .CDN(n3386), 
        .Q(serial_data_staging_1[11]) );
  dfcrq1 \serial_data_staging_1_reg[12]  ( .D(n2657), .CP(wb_clk_i), .CDN(
        n3379), .Q(serial_data_staging_1[12]) );
  dfcrq1 \serial_data_staging_2_reg[0]  ( .D(n2642), .CP(n3334), .CDN(n3386), 
        .Q(serial_data_staging_2[0]) );
  dfcrq1 \serial_data_staging_2_reg[1]  ( .D(n2641), .CP(wb_clk_i), .CDN(n3369), .Q(serial_data_staging_2[1]) );
  dfcrq1 \serial_data_staging_2_reg[2]  ( .D(n2640), .CP(n3334), .CDN(n3380), 
        .Q(serial_data_staging_2[2]) );
  dfcrq1 \serial_data_staging_2_reg[3]  ( .D(n2639), .CP(n3333), .CDN(n3348), 
        .Q(serial_data_staging_2[3]) );
  dfcrq1 \serial_data_staging_2_reg[4]  ( .D(n2638), .CP(n3334), .CDN(n3371), 
        .Q(serial_data_staging_2[4]) );
  dfcrq1 \serial_data_staging_2_reg[5]  ( .D(n2637), .CP(n3334), .CDN(n3376), 
        .Q(serial_data_staging_2[5]) );
  dfcrq1 \serial_data_staging_2_reg[6]  ( .D(n2636), .CP(n3332), .CDN(n3375), 
        .Q(serial_data_staging_2[6]) );
  dfcrq1 \serial_data_staging_2_reg[7]  ( .D(n2635), .CP(n3334), .CDN(n3338), 
        .Q(serial_data_staging_2[7]) );
  dfcrq1 \serial_data_staging_2_reg[8]  ( .D(n2634), .CP(n3334), .CDN(n3375), 
        .Q(serial_data_staging_2[8]) );
  dfcrq1 \serial_data_staging_2_reg[9]  ( .D(n2633), .CP(n3334), .CDN(n3346), 
        .Q(serial_data_staging_2[9]) );
  dfcrq1 \serial_data_staging_2_reg[10]  ( .D(n2632), .CP(n3334), .CDN(n3355), 
        .Q(serial_data_staging_2[10]) );
  dfcrq1 \serial_data_staging_2_reg[11]  ( .D(n2631), .CP(n3334), .CDN(n3387), 
        .Q(serial_data_staging_2[11]) );
  dfcrq1 \serial_data_staging_2_reg[12]  ( .D(n2630), .CP(n3334), .CDN(n3378), 
        .Q(serial_data_staging_2[12]) );
  dfcrq1 \pwr_ctrl_out_reg[0]  ( .D(n2600), .CP(n3298), .CDN(n3339), .Q(n432)
         );
  dfcrq1 \pwr_ctrl_out_reg[3]  ( .D(n2599), .CP(n3313), .CDN(n3378), .Q(n429)
         );
  dfcrq1 \pwr_ctrl_out_reg[2]  ( .D(n2598), .CP(n3299), .CDN(n3375), .Q(n430)
         );
  dfcrq1 \pwr_ctrl_out_reg[1]  ( .D(n2597), .CP(n3315), .CDN(n3380), .Q(n431)
         );
  dfcrq1 \mgmt_gpio_data_buf_reg[0]  ( .D(n2596), .CP(n3317), .CDN(n3365), .Q(
        mgmt_gpio_data_buf[0]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[1]  ( .D(n2595), .CP(n3315), .CDN(n3383), .Q(
        mgmt_gpio_data_buf[1]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[2]  ( .D(n2594), .CP(n3312), .CDN(n3382), .Q(
        mgmt_gpio_data_buf[2]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[3]  ( .D(n2593), .CP(n3324), .CDN(n3382), .Q(
        mgmt_gpio_data_buf[3]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[4]  ( .D(n2592), .CP(n3324), .CDN(n3382), .Q(
        mgmt_gpio_data_buf[4]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[5]  ( .D(n2591), .CP(n3324), .CDN(n3337), .Q(
        mgmt_gpio_data_buf[5]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[6]  ( .D(n2590), .CP(n3321), .CDN(n3337), .Q(
        mgmt_gpio_data_buf[6]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[7]  ( .D(n2589), .CP(n3300), .CDN(n3384), .Q(
        mgmt_gpio_data_buf[7]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[8]  ( .D(n2580), .CP(n3324), .CDN(n3381), .Q(
        mgmt_gpio_data_buf[8]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[9]  ( .D(n2579), .CP(n3324), .CDN(n3380), .Q(
        mgmt_gpio_data_buf[9]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[10]  ( .D(n2578), .CP(n3324), .CDN(n3338), 
        .Q(mgmt_gpio_data_buf[10]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[11]  ( .D(n2577), .CP(n3324), .CDN(n3381), 
        .Q(mgmt_gpio_data_buf[11]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[12]  ( .D(n2576), .CP(n3324), .CDN(n3343), 
        .Q(mgmt_gpio_data_buf[12]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[13]  ( .D(n2575), .CP(n3324), .CDN(n3385), 
        .Q(mgmt_gpio_data_buf[13]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[14]  ( .D(n2574), .CP(n3300), .CDN(n3345), 
        .Q(mgmt_gpio_data_buf[14]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[15]  ( .D(n2573), .CP(n3321), .CDN(n3336), 
        .Q(mgmt_gpio_data_buf[15]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[16]  ( .D(n2564), .CP(n3324), .CDN(n3375), 
        .Q(mgmt_gpio_data_buf[16]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[17]  ( .D(n2563), .CP(n3321), .CDN(n3357), 
        .Q(mgmt_gpio_data_buf[17]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[18]  ( .D(n2562), .CP(n3321), .CDN(n3383), 
        .Q(mgmt_gpio_data_buf[18]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[19]  ( .D(n2561), .CP(n3299), .CDN(n3377), 
        .Q(mgmt_gpio_data_buf[19]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[20]  ( .D(n2560), .CP(n3299), .CDN(n3377), 
        .Q(mgmt_gpio_data_buf[20]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[21]  ( .D(n2559), .CP(n3299), .CDN(n3379), 
        .Q(mgmt_gpio_data_buf[21]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[22]  ( .D(n2558), .CP(n3299), .CDN(n3363), 
        .Q(mgmt_gpio_data_buf[22]) );
  dfcrq1 \mgmt_gpio_data_buf_reg[23]  ( .D(n2557), .CP(n3299), .CDN(n3384), 
        .Q(mgmt_gpio_data_buf[23]) );
  dfcrq1 \mgmt_gpio_data_reg[31]  ( .D(n3048), .CP(n3299), .CDN(n3385), .Q(
        mgmt_gpio_out[31]) );
  dfcrq1 \mgmt_gpio_data_reg[30]  ( .D(n3047), .CP(n3299), .CDN(n3377), .Q(
        mgmt_gpio_out[30]) );
  dfcrq1 \mgmt_gpio_data_reg[29]  ( .D(n3046), .CP(n3299), .CDN(n3338), .Q(
        mgmt_gpio_out[29]) );
  dfcrq1 \mgmt_gpio_data_reg[28]  ( .D(n3045), .CP(n3309), .CDN(n3385), .Q(
        mgmt_gpio_out[28]) );
  dfcrq1 \mgmt_gpio_data_reg[27]  ( .D(n3044), .CP(n3310), .CDN(n3345), .Q(
        mgmt_gpio_out[27]) );
  dfcrq1 \mgmt_gpio_data_reg[26]  ( .D(n3043), .CP(n3304), .CDN(n3345), .Q(
        mgmt_gpio_out[26]) );
  dfcrq1 \mgmt_gpio_data_reg[25]  ( .D(n3042), .CP(n3298), .CDN(n3347), .Q(
        mgmt_gpio_out[25]) );
  dfcrq1 \mgmt_gpio_data_reg[24]  ( .D(n3041), .CP(n3313), .CDN(n3345), .Q(
        mgmt_gpio_out[24]) );
  dfcrq1 \mgmt_gpio_data_reg[0]  ( .D(n2588), .CP(n3299), .CDN(n3347), .Q(
        mgmt_gpio_data_0) );
  dfcrq1 \mgmt_gpio_data_reg[1]  ( .D(n2587), .CP(n3315), .CDN(n3345), .Q(
        mgmt_gpio_data_1) );
  dfcrq1 \mgmt_gpio_data_reg[2]  ( .D(n2586), .CP(n3317), .CDN(n3347), .Q(
        mgmt_gpio_out[2]) );
  dfcrq1 \mgmt_gpio_data_reg[3]  ( .D(n2585), .CP(n3298), .CDN(n3378), .Q(
        mgmt_gpio_out[3]) );
  dfcrq1 \mgmt_gpio_data_reg[4]  ( .D(n2584), .CP(n3298), .CDN(n3347), .Q(
        mgmt_gpio_out[4]) );
  dfcrq1 \mgmt_gpio_data_reg[5]  ( .D(n2583), .CP(n3298), .CDN(n3345), .Q(
        mgmt_gpio_out[5]) );
  dfcrq1 \mgmt_gpio_data_reg[6]  ( .D(n2582), .CP(n3298), .CDN(n3345), .Q(
        mgmt_gpio_data_6) );
  dfcrq1 \mgmt_gpio_data_reg[7]  ( .D(n2581), .CP(n3298), .CDN(n3380), .Q(
        mgmt_gpio_out[7]) );
  dfcrq1 \mgmt_gpio_data_reg[8]  ( .D(n2572), .CP(n3298), .CDN(n3337), .Q(
        mgmt_gpio_data_8) );
  dfcrq1 \mgmt_gpio_data_reg[9]  ( .D(n2571), .CP(n3298), .CDN(n3345), .Q(
        mgmt_gpio_data_9) );
  dfcrq1 \mgmt_gpio_data_reg[10]  ( .D(n2570), .CP(n3298), .CDN(n3347), .Q(
        mgmt_gpio_data_10) );
  dfcrq1 \mgmt_gpio_data_reg[11]  ( .D(n2569), .CP(n3298), .CDN(n3346), .Q(
        mgmt_gpio_out[11]) );
  dfcrq1 \mgmt_gpio_data_reg[12]  ( .D(n2568), .CP(n3303), .CDN(n3336), .Q(
        mgmt_gpio_out[12]) );
  dfcrq1 \mgmt_gpio_data_reg[13]  ( .D(n2567), .CP(n3315), .CDN(n3346), .Q(
        mgmt_gpio_data_13) );
  dfcrq1 \mgmt_gpio_data_reg[14]  ( .D(n2566), .CP(n3312), .CDN(n3368), .Q(
        mgmt_gpio_data_14) );
  dfcrq1 \mgmt_gpio_data_reg[15]  ( .D(n2565), .CP(n3313), .CDN(n3346), .Q(
        mgmt_gpio_data_15) );
  dfcrq1 \mgmt_gpio_data_reg[16]  ( .D(n2556), .CP(n3323), .CDN(n3347), .Q(
        mgmt_gpio_out[16]) );
  dfcrq1 \mgmt_gpio_data_reg[17]  ( .D(n2555), .CP(n3325), .CDN(n3346), .Q(
        mgmt_gpio_out[17]) );
  dfcrq1 \mgmt_gpio_data_reg[18]  ( .D(n2554), .CP(n3329), .CDN(n3347), .Q(
        mgmt_gpio_out[18]) );
  dfcrq1 \mgmt_gpio_data_reg[19]  ( .D(n2553), .CP(n3328), .CDN(n3346), .Q(
        mgmt_gpio_out[19]) );
  dfcrq1 \mgmt_gpio_data_reg[20]  ( .D(n2552), .CP(n3307), .CDN(n3346), .Q(
        mgmt_gpio_out[20]) );
  dfcrq1 \mgmt_gpio_data_reg[21]  ( .D(n2551), .CP(n3327), .CDN(n3357), .Q(
        mgmt_gpio_out[21]) );
  dfcrq1 \mgmt_gpio_data_reg[22]  ( .D(n2550), .CP(n3314), .CDN(n3347), .Q(
        mgmt_gpio_out[22]) );
  dfcrq1 \mgmt_gpio_data_reg[23]  ( .D(n2549), .CP(n3319), .CDN(n3346), .Q(
        mgmt_gpio_out[23]) );
  dfcrq1 \hkspi/pass_thru_mgmt_delay_reg  ( .D(n2534), .CP(n3291), .CDN(n3293), 
        .Q(pass_thru_mgmt_delay) );
  dfcrq1 \hkspi/pass_thru_user_delay_reg  ( .D(n2533), .CP(n3291), .CDN(n2523), 
        .Q(pass_thru_user_delay) );
  dfcrq1 \hkspi/writemode_reg  ( .D(n2532), .CP(n3291), .CDN(n3295), .Q(
        \hkspi/writemode ) );
  dfcrq1 \hkspi/predata_reg[0]  ( .D(n2531), .CP(n3291), .CDN(n2523), .Q(
        idata[1]) );
  dfcrq1 \hkspi/predata_reg[1]  ( .D(n2530), .CP(n3291), .CDN(n3295), .Q(
        idata[2]) );
  dfcrq1 \hkspi/predata_reg[2]  ( .D(n2529), .CP(n3291), .CDN(n2523), .Q(
        idata[3]) );
  dfcrq1 \hkspi/predata_reg[3]  ( .D(n2528), .CP(n3291), .CDN(n3294), .Q(
        idata[4]) );
  dfcrq1 \hkspi/predata_reg[4]  ( .D(n2527), .CP(n3291), .CDN(n3293), .Q(
        idata[5]) );
  dfcrq1 \hkspi/predata_reg[5]  ( .D(n2526), .CP(mgmt_gpio_in[4]), .CDN(n3295), 
        .Q(idata[6]) );
  dfcrq1 \hkspi/predata_reg[6]  ( .D(n2525), .CP(mgmt_gpio_in[4]), .CDN(n2523), 
        .Q(idata[7]) );
  dfcrq1 \hkspi/readmode_reg  ( .D(n2524), .CP(mgmt_gpio_in[4]), .CDN(n2523), 
        .Q(\hkspi/readmode ) );
  dfpfb1 \hkspi/sdoenb_reg  ( .D(\hkspi/N34 ), .CPN(n3291), .SDN(n3295), .Q(
        sdo_enb) );
  dfcfq1 \hkspi/wrstb_reg  ( .D(n3081), .CPN(mgmt_gpio_in[4]), .CDN(n2523), 
        .Q(wrstb) );
  dfcfq1 \hkspi/ldata_reg[0]  ( .D(n2548), .CPN(mgmt_gpio_in[4]), .CDN(n2523), 
        .Q(\hkspi/ldata[0] ) );
  dfcfq1 \hkspi/ldata_reg[1]  ( .D(n2547), .CPN(mgmt_gpio_in[4]), .CDN(n3295), 
        .Q(\hkspi/ldata[1] ) );
  dfcfq1 \hkspi/ldata_reg[2]  ( .D(n2546), .CPN(n3291), .CDN(n2523), .Q(
        \hkspi/ldata[2] ) );
  dfcfq1 \hkspi/ldata_reg[3]  ( .D(n2545), .CPN(n3291), .CDN(n2523), .Q(
        \hkspi/ldata[3] ) );
  dfcfq1 \hkspi/ldata_reg[4]  ( .D(n2544), .CPN(mgmt_gpio_in[4]), .CDN(n3295), 
        .Q(\hkspi/ldata[4] ) );
  dfcfq1 \hkspi/ldata_reg[5]  ( .D(n2543), .CPN(mgmt_gpio_in[4]), .CDN(n3295), 
        .Q(\hkspi/ldata[5] ) );
  dfcfq1 \hkspi/ldata_reg[6]  ( .D(n2542), .CPN(mgmt_gpio_in[4]), .CDN(n3295), 
        .Q(\hkspi/ldata[6] ) );
  dfcfq1 \hkspi/ldata_reg[7]  ( .D(n2541), .CPN(mgmt_gpio_in[4]), .CDN(n2523), 
        .Q(sdo) );
  dfcrn1 \gpio_configure_reg[4][10]  ( .D(n2522), .CP(n3310), .CDN(n3345), 
        .QN(\gpio_configure[4][10] ) );
  dfcrn1 \gpio_configure_reg[16][10]  ( .D(n2521), .CP(n3298), .CDN(n3347), 
        .QN(\gpio_configure[16][10] ) );
  dfcrn1 \gpio_configure_reg[15][1]  ( .D(n2520), .CP(n3299), .CDN(n3347), 
        .QN(\gpio_configure[15][1] ) );
  dfcrn1 \gpio_configure_reg[15][0]  ( .D(n2519), .CP(n3323), .CDN(n3346), 
        .QN(\gpio_configure[15][0] ) );
  dfcrn1 \gpio_configure_reg[0][12]  ( .D(n2518), .CP(n3318), .CDN(n3363), 
        .QN(\gpio_configure[0][12] ) );
  dfcrn1 \gpio_configure_reg[0][11]  ( .D(n2517), .CP(n3308), .CDN(n3346), 
        .QN(\gpio_configure[0][11] ) );
  dfcrn1 \gpio_configure_reg[8][10]  ( .D(n2516), .CP(n3309), .CDN(n3370), 
        .QN(\gpio_configure[8][10] ) );
  dfcrn1 \gpio_configure_reg[7][1]  ( .D(n2515), .CP(n3310), .CDN(n3346), .QN(
        \gpio_configure[7][1] ) );
  dfcrn1 \gpio_configure_reg[7][0]  ( .D(n2514), .CP(n3298), .CDN(n3355), .QN(
        \gpio_configure[7][0] ) );
  dfcrn1 \pll_trim_reg[7]  ( .D(n2513), .CP(n3299), .CDN(n3384), .QN(
        pll_trim[7]) );
  dfcrn1 \pll_trim_reg[6]  ( .D(n2512), .CP(n3315), .CDN(n3347), .QN(
        pll_trim[6]) );
  dfcrn1 \pll_trim_reg[5]  ( .D(n2511), .CP(n3301), .CDN(n3382), .QN(
        pll_trim[5]) );
  dfcrn1 \pll_trim_reg[4]  ( .D(n2510), .CP(n3324), .CDN(n3383), .QN(
        pll_trim[4]) );
  dfcrn1 \pll_trim_reg[3]  ( .D(n2509), .CP(n3304), .CDN(n3349), .QN(
        pll_trim[3]) );
  dfcrn1 \pll_trim_reg[2]  ( .D(n2508), .CP(n3322), .CDN(n3358), .QN(
        pll_trim[2]) );
  dfcrn1 \pll_trim_reg[1]  ( .D(n2507), .CP(n3329), .CDN(n3346), .QN(
        pll_trim[1]) );
  dfcrn1 \pll_trim_reg[0]  ( .D(n2506), .CP(n3316), .CDN(n3371), .QN(
        pll_trim[0]) );
  dfcrn1 \gpio_configure_reg[12][10]  ( .D(n2505), .CP(n3302), .CDN(n3346), 
        .QN(\gpio_configure[12][10] ) );
  dfcrn1 \gpio_configure_reg[11][1]  ( .D(n2504), .CP(n3301), .CDN(n3381), 
        .QN(\gpio_configure[11][1] ) );
  dfcrn1 \gpio_configure_reg[11][0]  ( .D(n2503), .CP(n3301), .CDN(n3364), 
        .QN(\gpio_configure[11][0] ) );
  dfcrn1 \gpio_configure_reg[36][12]  ( .D(n2502), .CP(n3318), .CDN(n3346), 
        .QN(\gpio_configure[36][12] ) );
  dfcrn1 \gpio_configure_reg[36][11]  ( .D(n2501), .CP(n3313), .CDN(n3369), 
        .QN(\gpio_configure[36][11] ) );
  dfcrn1 \gpio_configure_reg[35][1]  ( .D(n2500), .CP(n3302), .CDN(n3379), 
        .QN(\gpio_configure[35][1] ) );
  dfcrn1 \gpio_configure_reg[35][0]  ( .D(n2499), .CP(n3322), .CDN(n3345), 
        .QN(\gpio_configure[35][0] ) );
  dfcrn1 \gpio_configure_reg[20][10]  ( .D(n2498), .CP(csclk), .CDN(n3387), 
        .QN(\gpio_configure[20][10] ) );
  dfcrn1 \gpio_configure_reg[19][1]  ( .D(n2497), .CP(n3316), .CDN(n3347), 
        .QN(\gpio_configure[19][1] ) );
  dfcrn1 \gpio_configure_reg[19][0]  ( .D(n2496), .CP(n3316), .CDN(n3345), 
        .QN(\gpio_configure[19][0] ) );
  dfcrn1 \gpio_configure_reg[24][10]  ( .D(n2495), .CP(n3301), .CDN(n3345), 
        .QN(\gpio_configure[24][10] ) );
  dfcrn1 \gpio_configure_reg[23][1]  ( .D(n2494), .CP(n3308), .CDN(n3351), 
        .QN(\gpio_configure[23][1] ) );
  dfcrn1 \gpio_configure_reg[23][0]  ( .D(n2493), .CP(n3301), .CDN(n3366), 
        .QN(\gpio_configure[23][0] ) );
  dfcrn1 \gpio_configure_reg[32][10]  ( .D(n2492), .CP(n3322), .CDN(n3350), 
        .QN(\gpio_configure[32][10] ) );
  dfcrn1 \gpio_configure_reg[31][1]  ( .D(n2491), .CP(n3302), .CDN(n3365), 
        .QN(\gpio_configure[31][1] ) );
  dfcrn1 \gpio_configure_reg[31][0]  ( .D(n2490), .CP(n3322), .CDN(n3345), 
        .QN(\gpio_configure[31][0] ) );
  dfcrn1 \gpio_configure_reg[28][10]  ( .D(n2489), .CP(n3315), .CDN(n3347), 
        .QN(\gpio_configure[28][10] ) );
  dfcrn1 \gpio_configure_reg[27][1]  ( .D(n2488), .CP(n3316), .CDN(n3386), 
        .QN(\gpio_configure[27][1] ) );
  dfcrn1 \gpio_configure_reg[27][0]  ( .D(n2487), .CP(n3329), .CDN(n3345), 
        .QN(\gpio_configure[27][0] ) );
  dfcrn1 \pad_count_2_reg[0]  ( .D(n2540), .CP(n3332), .CDN(n3377), .QN(
        pad_count_2[0]) );
  dfcrn1 \pad_count_2_reg[1]  ( .D(n2539), .CP(n3332), .CDN(n3348), .QN(
        pad_count_2[1]) );
  dfcrn1 \pad_count_2_reg[4]  ( .D(n2538), .CP(n3332), .CDN(n3376), .QN(
        pad_count_2[4]) );
  dfcrn1 \pad_count_1_reg[1]  ( .D(n2537), .CP(n3332), .CDN(n3356), .QN(
        pad_count_1[1]) );
  dfcrn1 \pad_count_1_reg[4]  ( .D(n2536), .CP(n3332), .CDN(n3347), .QN(
        pad_count_1[4]) );
  dfcrn1 \gpio_configure_reg[11][10]  ( .D(n2486), .CP(n3314), .CDN(n3385), 
        .QN(\gpio_configure[11][10] ) );
  dfcrn1 \gpio_configure_reg[10][1]  ( .D(n2485), .CP(n3299), .CDN(n473), .QN(
        \gpio_configure[10][1] ) );
  dfcrn1 \gpio_configure_reg[10][0]  ( .D(n2484), .CP(n3306), .CDN(n474), .QN(
        \gpio_configure[10][0] ) );
  dfcrn1 \pll_div_reg[2]  ( .D(n2483), .CP(n3298), .CDN(n3344), .QN(pll_div[2]) );
  dfcrn1 \gpio_configure_reg[3][11]  ( .D(n2482), .CP(n3309), .CDN(n473), .QN(
        \gpio_configure[3][11] ) );
  dfcrn1 \gpio_configure_reg[7][10]  ( .D(n2481), .CP(n3323), .CDN(n474), .QN(
        \gpio_configure[7][10] ) );
  dfcrn1 \gpio_configure_reg[6][1]  ( .D(n2480), .CP(n3319), .CDN(n3344), .QN(
        \gpio_configure[6][1] ) );
  dfcrn1 \gpio_configure_reg[6][0]  ( .D(n2479), .CP(n3322), .CDN(n473), .QN(
        \gpio_configure[6][0] ) );
  dfcrn1 \gpio_configure_reg[15][10]  ( .D(n2478), .CP(n3322), .CDN(n474), 
        .QN(\gpio_configure[15][10] ) );
  dfcrn1 \gpio_configure_reg[14][1]  ( .D(n2477), .CP(n3316), .CDN(n3344), 
        .QN(\gpio_configure[14][1] ) );
  dfcrn1 \gpio_configure_reg[14][0]  ( .D(n2476), .CP(n3302), .CDN(n3343), 
        .QN(\gpio_configure[14][0] ) );
  dfcrn1 \gpio_configure_reg[35][10]  ( .D(n2475), .CP(n3301), .CDN(n3343), 
        .QN(\gpio_configure[35][10] ) );
  dfcrn1 \gpio_configure_reg[34][1]  ( .D(n2474), .CP(n3300), .CDN(n3342), 
        .QN(\gpio_configure[34][1] ) );
  dfcrn1 \gpio_configure_reg[34][0]  ( .D(n2473), .CP(n3329), .CDN(n3341), 
        .QN(\gpio_configure[34][0] ) );
  dfcrn1 \gpio_configure_reg[19][10]  ( .D(n2472), .CP(n3322), .CDN(n473), 
        .QN(\gpio_configure[19][10] ) );
  dfcrn1 \gpio_configure_reg[18][1]  ( .D(n2471), .CP(n3322), .CDN(n3342), 
        .QN(\gpio_configure[18][1] ) );
  dfcrn1 \gpio_configure_reg[18][0]  ( .D(n2470), .CP(n3322), .CDN(n3341), 
        .QN(\gpio_configure[18][0] ) );
  dfcrn1 \gpio_configure_reg[23][10]  ( .D(n2469), .CP(n3322), .CDN(n3344), 
        .QN(\gpio_configure[23][10] ) );
  dfcrn1 \gpio_configure_reg[22][1]  ( .D(n2468), .CP(n3322), .CDN(n3343), 
        .QN(\gpio_configure[22][1] ) );
  dfcrn1 \gpio_configure_reg[22][0]  ( .D(n2467), .CP(n3322), .CDN(n3340), 
        .QN(\gpio_configure[22][0] ) );
  dfcrn1 \gpio_configure_reg[31][10]  ( .D(n2466), .CP(n3304), .CDN(n3340), 
        .QN(\gpio_configure[31][10] ) );
  dfcrn1 \gpio_configure_reg[30][1]  ( .D(n2465), .CP(n3316), .CDN(n3340), 
        .QN(\gpio_configure[30][1] ) );
  dfcrn1 \gpio_configure_reg[30][0]  ( .D(n2464), .CP(n3302), .CDN(n3340), 
        .QN(\gpio_configure[30][0] ) );
  dfcrn1 \gpio_configure_reg[27][10]  ( .D(n2463), .CP(n3297), .CDN(n3340), 
        .QN(\gpio_configure[27][10] ) );
  dfcrn1 \gpio_configure_reg[26][1]  ( .D(n2462), .CP(n3297), .CDN(n3340), 
        .QN(\gpio_configure[26][1] ) );
  dfcrn1 \gpio_configure_reg[26][0]  ( .D(n2461), .CP(n3297), .CDN(n3340), 
        .QN(\gpio_configure[26][0] ) );
  dfcrn1 \gpio_configure_reg[14][10]  ( .D(n2460), .CP(n3297), .CDN(n3342), 
        .QN(\gpio_configure[14][10] ) );
  dfcrn1 \gpio_configure_reg[13][1]  ( .D(n2459), .CP(n3297), .CDN(n3341), 
        .QN(\gpio_configure[13][1] ) );
  dfcrn1 \gpio_configure_reg[13][0]  ( .D(n2458), .CP(n3297), .CDN(n474), .QN(
        \gpio_configure[13][0] ) );
  dfcrn1 \gpio_configure_reg[10][10]  ( .D(n2457), .CP(n3297), .CDN(n3340), 
        .QN(\gpio_configure[10][10] ) );
  dfcrn1 \gpio_configure_reg[9][1]  ( .D(n2456), .CP(n3297), .CDN(n3343), .QN(
        \gpio_configure[9][1] ) );
  dfcrn1 \gpio_configure_reg[9][0]  ( .D(n2455), .CP(n3313), .CDN(n3342), .QN(
        \gpio_configure[9][0] ) );
  dfcrn1 \pll_trim_reg[25]  ( .D(n2454), .CP(n3299), .CDN(n3341), .QN(
        pll_trim[25]) );
  dfcrn1 \pll_trim_reg[24]  ( .D(n2453), .CP(n3321), .CDN(n473), .QN(
        pll_trim[24]) );
  dfcrn1 \pll_sel_reg[1]  ( .D(n2452), .CP(n3324), .CDN(n3340), .QN(pll_sel[1]) );
  dfcrn1 \pll90_sel_reg[1]  ( .D(n2451), .CP(n3300), .CDN(n3343), .QN(
        pll90_sel[1]) );
  dfcrn1 \gpio_configure_reg[6][10]  ( .D(n2450), .CP(n3297), .CDN(n3342), 
        .QN(\gpio_configure[6][10] ) );
  dfcrn1 \gpio_configure_reg[5][1]  ( .D(n2449), .CP(n3312), .CDN(n3341), .QN(
        \gpio_configure[5][1] ) );
  dfcrn1 \gpio_configure_reg[5][0]  ( .D(n2448), .CP(n3298), .CDN(n3344), .QN(
        \gpio_configure[5][0] ) );
  dfcrn1 pll_dco_ena_reg ( .D(n2447), .CP(n3321), .CDN(n3340), .QN(pll_dco_ena) );
  dfcrn1 pll_bypass_reg ( .D(n2446), .CP(n3297), .CDN(n3343), .QN(pll_bypass)
         );
  dfcrn1 \gpio_configure_reg[2][10]  ( .D(n2445), .CP(n3300), .CDN(n3342), 
        .QN(\gpio_configure[2][10] ) );
  dfcrn1 \gpio_configure_reg[37][1]  ( .D(n2444), .CP(n3321), .CDN(n3341), 
        .QN(\gpio_configure[37][1] ) );
  dfcrn1 \gpio_configure_reg[37][0]  ( .D(n2443), .CP(n3297), .CDN(n474), .QN(
        \gpio_configure[37][0] ) );
  dfcrn1 \gpio_configure_reg[22][10]  ( .D(n2442), .CP(n3297), .CDN(n3340), 
        .QN(\gpio_configure[22][10] ) );
  dfcrn1 \gpio_configure_reg[21][1]  ( .D(n2441), .CP(n3320), .CDN(n3343), 
        .QN(\gpio_configure[21][1] ) );
  dfcrn1 \gpio_configure_reg[21][0]  ( .D(n2440), .CP(n3321), .CDN(n3342), 
        .QN(\gpio_configure[21][0] ) );
  dfcrn1 \gpio_configure_reg[34][10]  ( .D(n2439), .CP(csclk), .CDN(n3341), 
        .QN(\gpio_configure[34][10] ) );
  dfcrn1 \gpio_configure_reg[33][1]  ( .D(n2438), .CP(csclk), .CDN(n3344), 
        .QN(\gpio_configure[33][1] ) );
  dfcrn1 \gpio_configure_reg[33][0]  ( .D(n2437), .CP(csclk), .CDN(n3340), 
        .QN(\gpio_configure[33][0] ) );
  dfcrn1 \gpio_configure_reg[18][10]  ( .D(n2436), .CP(csclk), .CDN(n3343), 
        .QN(\gpio_configure[18][10] ) );
  dfcrn1 \gpio_configure_reg[17][1]  ( .D(n2435), .CP(csclk), .CDN(n3342), 
        .QN(\gpio_configure[17][1] ) );
  dfcrn1 \gpio_configure_reg[17][0]  ( .D(n2434), .CP(n3301), .CDN(n3341), 
        .QN(\gpio_configure[17][0] ) );
  dfcrn1 \gpio_configure_reg[30][10]  ( .D(n2433), .CP(n3301), .CDN(n474), 
        .QN(\gpio_configure[30][10] ) );
  dfcrn1 \gpio_configure_reg[29][1]  ( .D(n2432), .CP(n3302), .CDN(n3340), 
        .QN(\gpio_configure[29][1] ) );
  dfcrn1 \gpio_configure_reg[29][0]  ( .D(n2431), .CP(n3297), .CDN(n3343), 
        .QN(\gpio_configure[29][0] ) );
  dfcrn1 \gpio_configure_reg[26][10]  ( .D(n2430), .CP(n3320), .CDN(n3342), 
        .QN(\gpio_configure[26][10] ) );
  dfcrn1 \gpio_configure_reg[25][1]  ( .D(n2429), .CP(n3321), .CDN(n3341), 
        .QN(\gpio_configure[25][1] ) );
  dfcrn1 \gpio_configure_reg[25][0]  ( .D(n2428), .CP(n3303), .CDN(n473), .QN(
        \gpio_configure[25][0] ) );
  dfcrn1 \gpio_configure_reg[5][10]  ( .D(n2427), .CP(n3297), .CDN(n3340), 
        .QN(\gpio_configure[5][10] ) );
  dfcrn1 \gpio_configure_reg[4][1]  ( .D(n2426), .CP(n3321), .CDN(n3343), .QN(
        \gpio_configure[4][1] ) );
  dfcrn1 \gpio_configure_reg[4][0]  ( .D(n2425), .CP(n3297), .CDN(porb), .QN(
        \gpio_configure[4][0] ) );
  dfcrn1 \gpio_configure_reg[13][10]  ( .D(n2424), .CP(n3312), .CDN(porb), 
        .QN(\gpio_configure[13][10] ) );
  dfcrn1 \gpio_configure_reg[12][1]  ( .D(n2423), .CP(n3303), .CDN(porb), .QN(
        \gpio_configure[12][1] ) );
  dfcrn1 \gpio_configure_reg[12][0]  ( .D(n2422), .CP(n3297), .CDN(porb), .QN(
        \gpio_configure[12][0] ) );
  dfcrn1 \gpio_configure_reg[17][10]  ( .D(n2421), .CP(n3297), .CDN(porb), 
        .QN(\gpio_configure[17][10] ) );
  dfcrn1 \gpio_configure_reg[16][1]  ( .D(n2420), .CP(n3320), .CDN(porb), .QN(
        \gpio_configure[16][1] ) );
  dfcrn1 \gpio_configure_reg[16][0]  ( .D(n2419), .CP(n3297), .CDN(porb), .QN(
        \gpio_configure[16][0] ) );
  dfcrn1 \gpio_configure_reg[1][12]  ( .D(n2418), .CP(n3321), .CDN(porb), .QN(
        \gpio_configure[1][12] ) );
  dfcrn1 \gpio_configure_reg[1][11]  ( .D(n2417), .CP(n3299), .CDN(porb), .QN(
        \gpio_configure[1][11] ) );
  dfcrn1 \gpio_configure_reg[0][1]  ( .D(n2416), .CP(n3321), .CDN(porb), .QN(
        \gpio_configure[0][1] ) );
  dfcrn1 \gpio_configure_reg[0][0]  ( .D(n2415), .CP(n3320), .CDN(n3338), .QN(
        \gpio_configure[0][0] ) );
  dfcrn1 \gpio_configure_reg[9][10]  ( .D(n2414), .CP(n3317), .CDN(n3339), 
        .QN(\gpio_configure[9][10] ) );
  dfcrn1 \gpio_configure_reg[8][1]  ( .D(n2413), .CP(n3320), .CDN(n3337), .QN(
        \gpio_configure[8][1] ) );
  dfcrn1 \gpio_configure_reg[8][0]  ( .D(n2412), .CP(n3303), .CDN(n3336), .QN(
        \gpio_configure[8][0] ) );
  dfcrn1 \pll_trim_reg[23]  ( .D(n2411), .CP(n3317), .CDN(n3338), .QN(
        pll_trim[23]) );
  dfcrn1 \pll_trim_reg[22]  ( .D(n2410), .CP(n3315), .CDN(n3339), .QN(
        pll_trim[22]) );
  dfcrn1 \pll_trim_reg[21]  ( .D(n2409), .CP(n3312), .CDN(n3337), .QN(
        pll_trim[21]) );
  dfcrn1 \pll_trim_reg[20]  ( .D(n2408), .CP(n3313), .CDN(n3336), .QN(
        pll_trim[20]) );
  dfcrn1 \pll_trim_reg[19]  ( .D(n2407), .CP(n3320), .CDN(n3338), .QN(
        pll_trim[19]) );
  dfcrn1 \pll_trim_reg[18]  ( .D(n2406), .CP(n3320), .CDN(n3339), .QN(
        pll_trim[18]) );
  dfcrn1 \pll_trim_reg[17]  ( .D(n2405), .CP(n3320), .CDN(n3337), .QN(
        pll_trim[17]) );
  dfcrn1 \pll_trim_reg[16]  ( .D(n2404), .CP(n3320), .CDN(n3336), .QN(
        pll_trim[16]) );
  dfcrn1 \pll_trim_reg[15]  ( .D(n2403), .CP(n3320), .CDN(n3338), .QN(
        pll_trim[15]) );
  dfcrn1 \pll_trim_reg[14]  ( .D(n2402), .CP(n3303), .CDN(n3339), .QN(
        pll_trim[14]) );
  dfcrn1 \pll_trim_reg[13]  ( .D(n2401), .CP(n3317), .CDN(n3337), .QN(
        pll_trim[13]) );
  dfcrn1 \pll_trim_reg[11]  ( .D(n2400), .CP(n3315), .CDN(n3336), .QN(
        pll_trim[11]) );
  dfcrn1 \pll_trim_reg[10]  ( .D(n2399), .CP(n3314), .CDN(n3338), .QN(
        pll_trim[10]) );
  dfcrn1 \pll_trim_reg[9]  ( .D(n2398), .CP(n3316), .CDN(n3339), .QN(
        pll_trim[9]) );
  dfcrn1 \pll_trim_reg[8]  ( .D(n2397), .CP(n3301), .CDN(n3337), .QN(
        pll_trim[8]) );
  dfcrn1 \gpio_configure_reg[25][10]  ( .D(n2396), .CP(n3302), .CDN(n3336), 
        .QN(\gpio_configure[25][10] ) );
  dfcrn1 \gpio_configure_reg[24][1]  ( .D(n2395), .CP(n3322), .CDN(n3379), 
        .QN(\gpio_configure[24][1] ) );
  dfcrn1 \gpio_configure_reg[24][0]  ( .D(n2394), .CP(n3320), .CDN(n3379), 
        .QN(\gpio_configure[24][0] ) );
  dfcrn1 \gpio_configure_reg[37][12]  ( .D(n2393), .CP(n3303), .CDN(n3379), 
        .QN(\gpio_configure[37][12] ) );
  dfcrn1 \gpio_configure_reg[37][11]  ( .D(n2392), .CP(n3325), .CDN(n3379), 
        .QN(\gpio_configure[37][11] ) );
  dfcrn1 \gpio_configure_reg[36][1]  ( .D(n2391), .CP(n3320), .CDN(n3379), 
        .QN(\gpio_configure[36][1] ) );
  dfcrn1 \gpio_configure_reg[36][0]  ( .D(n2390), .CP(n3312), .CDN(n3379), 
        .QN(\gpio_configure[36][0] ) );
  dfcrn1 \gpio_configure_reg[21][10]  ( .D(n2389), .CP(n3317), .CDN(n3379), 
        .QN(\gpio_configure[21][10] ) );
  dfcrn1 \gpio_configure_reg[20][1]  ( .D(n2388), .CP(n3315), .CDN(n3379), 
        .QN(\gpio_configure[20][1] ) );
  dfcrn1 \gpio_configure_reg[20][0]  ( .D(n2387), .CP(n3312), .CDN(n3379), 
        .QN(\gpio_configure[20][0] ) );
  dfcrn1 \gpio_configure_reg[33][10]  ( .D(n2386), .CP(n3313), .CDN(n3379), 
        .QN(\gpio_configure[33][10] ) );
  dfcrn1 \gpio_configure_reg[32][1]  ( .D(n2385), .CP(n3303), .CDN(n3338), 
        .QN(\gpio_configure[32][1] ) );
  dfcrn1 \gpio_configure_reg[32][0]  ( .D(n2384), .CP(n3320), .CDN(n3339), 
        .QN(\gpio_configure[32][0] ) );
  dfcrn1 \gpio_configure_reg[29][10]  ( .D(n2383), .CP(n3322), .CDN(n3337), 
        .QN(\gpio_configure[29][10] ) );
  dfcrn1 \gpio_configure_reg[28][1]  ( .D(n2382), .CP(n3304), .CDN(n3336), 
        .QN(\gpio_configure[28][1] ) );
  dfcrn1 \gpio_configure_reg[28][0]  ( .D(n2381), .CP(n3313), .CDN(n3338), 
        .QN(\gpio_configure[28][0] ) );
  dfcrn1 \gpio_configure_reg[3][0]  ( .D(n2380), .CP(n3302), .CDN(n3339), .QN(
        \gpio_configure[3][0] ) );
  dfcrn1 \gpio_configure_reg[2][1]  ( .D(n2379), .CP(n3316), .CDN(n3337), .QN(
        \gpio_configure[2][1] ) );
  dfcrn1 \gpio_configure_reg[2][0]  ( .D(n2378), .CP(n3301), .CDN(n3336), .QN(
        \gpio_configure[2][0] ) );
  dfcrn1 \gpio_configure_reg[1][1]  ( .D(n2377), .CP(n3322), .CDN(n3338), .QN(
        \gpio_configure[1][1] ) );
  dfcrn1 \gpio_configure_reg[1][0]  ( .D(n2376), .CP(n3327), .CDN(n3339), .QN(
        \gpio_configure[1][0] ) );
  dfnrq1 \wb_dat_o_reg[7]  ( .D(n2375), .CP(n3332), .Q(wb_dat_o[7]) );
  dfnrq1 \wb_dat_o_reg[15]  ( .D(n2374), .CP(n3332), .Q(wb_dat_o[15]) );
  dfnrq1 \wb_dat_o_reg[23]  ( .D(n2373), .CP(n3332), .Q(wb_dat_o[23]) );
  dfnrq1 \wb_dat_o_reg[31]  ( .D(n2372), .CP(n3332), .Q(wb_dat_o[31]) );
  dfnrq1 \wb_dat_o_reg[4]  ( .D(n2371), .CP(n3332), .Q(wb_dat_o[4]) );
  dfnrq1 \wb_dat_o_reg[12]  ( .D(n2370), .CP(n3332), .Q(wb_dat_o[12]) );
  dfnrq1 \wb_dat_o_reg[20]  ( .D(n2369), .CP(n3332), .Q(wb_dat_o[20]) );
  dfnrq1 \wb_dat_o_reg[28]  ( .D(n2368), .CP(n3332), .Q(wb_dat_o[28]) );
  dfnrq1 \wb_dat_o_reg[5]  ( .D(n2367), .CP(n3333), .Q(wb_dat_o[5]) );
  dfnrq1 \wb_dat_o_reg[13]  ( .D(n2366), .CP(n3333), .Q(wb_dat_o[13]) );
  dfnrq1 \wb_dat_o_reg[21]  ( .D(n2365), .CP(n3333), .Q(wb_dat_o[21]) );
  dfnrq1 \wb_dat_o_reg[29]  ( .D(n2364), .CP(n3333), .Q(wb_dat_o[29]) );
  dfnrq1 \wb_dat_o_reg[6]  ( .D(n2363), .CP(n3333), .Q(wb_dat_o[6]) );
  dfnrq1 \wb_dat_o_reg[14]  ( .D(n2362), .CP(n3333), .Q(wb_dat_o[14]) );
  dfnrq1 \wb_dat_o_reg[22]  ( .D(n2361), .CP(n3333), .Q(wb_dat_o[22]) );
  dfnrq1 \wb_dat_o_reg[30]  ( .D(n2360), .CP(n3333), .Q(wb_dat_o[30]) );
  dfnrq1 \wb_dat_o_reg[0]  ( .D(n2359), .CP(n3333), .Q(wb_dat_o[0]) );
  dfnrq1 \wb_dat_o_reg[8]  ( .D(n2358), .CP(n3333), .Q(wb_dat_o[8]) );
  dfnrq1 \wb_dat_o_reg[16]  ( .D(n2357), .CP(n3333), .Q(wb_dat_o[16]) );
  dfnrq1 \wb_dat_o_reg[24]  ( .D(n2356), .CP(n3333), .Q(wb_dat_o[24]) );
  dfnrq1 \wb_dat_o_reg[3]  ( .D(n2355), .CP(n3333), .Q(wb_dat_o[3]) );
  dfnrq1 \wb_dat_o_reg[11]  ( .D(n2354), .CP(n3333), .Q(wb_dat_o[11]) );
  dfnrq1 \wb_dat_o_reg[19]  ( .D(n2353), .CP(n3333), .Q(wb_dat_o[19]) );
  dfnrq1 \wb_dat_o_reg[27]  ( .D(n2352), .CP(n3333), .Q(wb_dat_o[27]) );
  dfnrq1 \wb_dat_o_reg[2]  ( .D(n2351), .CP(n3334), .Q(wb_dat_o[2]) );
  dfnrq1 \wb_dat_o_reg[10]  ( .D(n2350), .CP(n3330), .Q(wb_dat_o[10]) );
  dfnrq1 \wb_dat_o_reg[18]  ( .D(n2349), .CP(n3331), .Q(wb_dat_o[18]) );
  dfnrq1 \wb_dat_o_reg[26]  ( .D(n2348), .CP(n3332), .Q(wb_dat_o[26]) );
  dfnrq1 \wb_dat_o_reg[1]  ( .D(n2347), .CP(n3331), .Q(wb_dat_o[1]) );
  dfnrq1 \wb_dat_o_reg[9]  ( .D(n2346), .CP(n3333), .Q(wb_dat_o[9]) );
  dfnrq1 \wb_dat_o_reg[17]  ( .D(n2345), .CP(n3334), .Q(wb_dat_o[17]) );
  dfnrq1 \wb_dat_o_reg[25]  ( .D(n2344), .CP(n3330), .Q(wb_dat_o[25]) );
  oaim22d1 U519 ( .A1(n633), .A2(n3296), .B1(n620), .B2(mgmt_gpio_in[12]), 
        .ZN(n386) );
  aoi22d1 U3105 ( .A1(pass_thru_user), .A2(n3296), .B1(n2319), .B2(n2335), 
        .ZN(mgmt_gpio_out_9_prebuff) );
  inv0d0 U3108 ( .I(wb_clk_i), .ZN(n2322) );
  oan211d1 U3138 ( .C1(n3296), .C2(n2342), .B(n2341), .A(n2340), .ZN(csclk) );
  dfcrq1 wbbd_busy_reg ( .D(n3060), .CP(wb_clk_i), .CDN(n3292), .Q(wbbd_busy)
         );
  mx02d1 U3139 ( .I0(serial_load_pre), .I1(serial_bb_load), .S(
        serial_bb_enable), .Z(serial_load) );
  mx02d1 U3140 ( .I0(1'b1), .I1(mgmt_gpio_in[3]), .S(spi_is_enabled), .Z(
        \_1_net_[0] ) );
  aoim22d1 U3 ( .A1(n3265), .A2(n1701), .B1(\gpio_configure[3][5] ), .B2(n3265), .Z(n2690) );
  aoim22d1 U4 ( .A1(n3198), .A2(n1701), .B1(\gpio_configure[17][5] ), .B2(
        n3198), .Z(n2830) );
  aoim22d1 U5 ( .A1(n3147), .A2(n1701), .B1(\gpio_configure[18][5] ), .B2(
        n3147), .Z(n2840) );
  aoim22d1 U6 ( .A1(n2332), .A2(n1701), .B1(\gpio_configure[7][5] ), .B2(n2332), .Z(n2730) );
  aoim22d1 U7 ( .A1(n3168), .A2(n1701), .B1(\gpio_configure[9][5] ), .B2(n3168), .Z(n2750) );
  aoim22d1 U8 ( .A1(n3219), .A2(n1701), .B1(\gpio_configure[16][5] ), .B2(
        n3219), .Z(n2820) );
  aoim22d1 U9 ( .A1(n2326), .A2(n1701), .B1(\gpio_configure[15][5] ), .B2(
        n2326), .Z(n2810) );
  aoim22d1 U10 ( .A1(n3135), .A2(n1701), .B1(\gpio_configure[6][5] ), .B2(
        n3135), .Z(n2720) );
  aoim22d1 U11 ( .A1(n3164), .A2(n1701), .B1(\gpio_configure[13][5] ), .B2(
        n3164), .Z(n2790) );
  aoim22d1 U12 ( .A1(n2535), .A2(n1701), .B1(\gpio_configure[11][5] ), .B2(
        n2535), .Z(n2770) );
  aoim22d1 U13 ( .A1(n3139), .A2(n1701), .B1(\gpio_configure[14][5] ), .B2(
        n3139), .Z(n2800) );
  aoim22d1 U14 ( .A1(n3215), .A2(n1701), .B1(\gpio_configure[12][5] ), .B2(
        n3215), .Z(n2780) );
  aoim22d1 U15 ( .A1(n3211), .A2(n1701), .B1(\gpio_configure[4][5] ), .B2(
        n3211), .Z(n2700) );
  aoim22d1 U16 ( .A1(n3127), .A2(n1701), .B1(\gpio_configure[10][5] ), .B2(
        n3127), .Z(n2760) );
  aoim22d1 U17 ( .A1(n3273), .A2(n1701), .B1(\gpio_configure[1][5] ), .B2(
        n3273), .Z(n2670) );
  aoim22d1 U18 ( .A1(n824), .A2(n1701), .B1(mgmt_gpio_data[37]), .B2(n824), 
        .Z(n3054) );
  aoim22d1 U19 ( .A1(n3174), .A2(n1701), .B1(pll90_sel[2]), .B2(n3174), .Z(
        n2613) );
  inv0d0 U20 ( .I(n1541), .ZN(n1642) );
  aoi22d1 U21 ( .A1(n2267), .A2(\gpio_configure[17][0] ), .B1(n858), .B2(
        pll_ena), .ZN(n1797) );
  inv0d4 U22 ( .I(n1696), .ZN(n1646) );
  clk2d2 U23 ( .CLK(n482), .CN(n473), .C(n472) );
  inv0d0 U24 ( .I(n472), .ZN(n474) );
  inv0d1 U25 ( .I(n1815), .ZN(n2267) );
  nd04d0 U26 ( .A1(n735), .A2(n734), .A3(n733), .A4(n732), .ZN(n752) );
  nd04d0 U27 ( .A1(n785), .A2(n625), .A3(n733), .A4(n676), .ZN(n763) );
  nd04d0 U28 ( .A1(N863), .A2(n766), .A3(n765), .A4(n764), .ZN(n772) );
  nd04d0 U29 ( .A1(n570), .A2(n569), .A3(n568), .A4(n567), .ZN(n571) );
  nd04d0 U30 ( .A1(n1948), .A2(n1947), .A3(n1946), .A4(n1945), .ZN(n1999) );
  nd04d0 U31 ( .A1(n2015), .A2(n2014), .A3(n2013), .A4(n2012), .ZN(n2065) );
  nd04d0 U32 ( .A1(n2086), .A2(n2085), .A3(n2084), .A4(n2083), .ZN(n2136) );
  nd04d0 U33 ( .A1(n2114), .A2(n2113), .A3(n2112), .A4(n2111), .ZN(n2130) );
  nd04d0 U34 ( .A1(n943), .A2(n942), .A3(n941), .A4(n940), .ZN(n959) );
  nd04d0 U35 ( .A1(n2146), .A2(n2145), .A3(n2144), .A4(n2143), .ZN(n2157) );
  nd04d0 U36 ( .A1(n922), .A2(n921), .A3(n920), .A4(n919), .ZN(n938) );
  nd04d0 U37 ( .A1(n2168), .A2(n2167), .A3(n2166), .A4(n2165), .ZN(n2169) );
  nd04d0 U38 ( .A1(n2199), .A2(n2198), .A3(n2197), .A4(n2196), .ZN(n2214) );
  nd04d0 U39 ( .A1(n2273), .A2(n2272), .A3(n2271), .A4(n2270), .ZN(n2274) );
  nd04d0 U40 ( .A1(n926), .A2(n925), .A3(n924), .A4(n923), .ZN(n937) );
  nd04d0 U41 ( .A1(n930), .A2(n929), .A3(n928), .A4(n927), .ZN(n936) );
  nd04d0 U42 ( .A1(n934), .A2(n933), .A3(n932), .A4(n931), .ZN(n935) );
  nd04d0 U43 ( .A1(n1429), .A2(n1428), .A3(n1427), .A4(n1426), .ZN(n1445) );
  nd04d0 U44 ( .A1(n1433), .A2(n1432), .A3(n1431), .A4(n1430), .ZN(n1444) );
  nd04d0 U45 ( .A1(n1375), .A2(n1374), .A3(n1373), .A4(n1372), .ZN(n1386) );
  nd04d0 U46 ( .A1(n1494), .A2(n1493), .A3(n1492), .A4(n1491), .ZN(n1505) );
  nd04d0 U47 ( .A1(n1471), .A2(n1470), .A3(n1469), .A4(n1468), .ZN(n1472) );
  nd04d0 U48 ( .A1(n1942), .A2(n1941), .A3(n1940), .A4(n1939), .ZN(n1943) );
  nd04d0 U49 ( .A1(n1322), .A2(n1321), .A3(n1320), .A4(n1319), .ZN(n1328) );
  nd04d0 U50 ( .A1(n1938), .A2(n1937), .A3(n1936), .A4(n1935), .ZN(n1944) );
  nd04d0 U51 ( .A1(n1960), .A2(n1959), .A3(n1958), .A4(n1957), .ZN(n1961) );
  nd04d0 U52 ( .A1(n1259), .A2(n1258), .A3(n1257), .A4(n1256), .ZN(n1275) );
  nd04d0 U53 ( .A1(n1379), .A2(n1378), .A3(n1377), .A4(n1376), .ZN(n1385) );
  nd04d0 U54 ( .A1(n1884), .A2(n1883), .A3(n1882), .A4(n1881), .ZN(n1890) );
  nd04d0 U55 ( .A1(n1871), .A2(n1870), .A3(n1869), .A4(n1868), .ZN(n1872) );
  nd04d0 U56 ( .A1(n1867), .A2(n1866), .A3(n1865), .A4(n1864), .ZN(n1873) );
  nd04d0 U57 ( .A1(n1820), .A2(n1819), .A3(n1818), .A4(n1817), .ZN(n1821) );
  nd04d0 U58 ( .A1(n1814), .A2(n1813), .A3(n1812), .A4(n1811), .ZN(n1822) );
  nd04d0 U59 ( .A1(n1563), .A2(n1562), .A3(n1561), .A4(n1560), .ZN(n1564) );
  nd04d0 U60 ( .A1(n1520), .A2(n1519), .A3(n1518), .A4(n1517), .ZN(n1536) );
  nd04d0 U61 ( .A1(n1850), .A2(n1849), .A3(n1848), .A4(n1847), .ZN(n1851) );
  nd04d0 U62 ( .A1(n1524), .A2(n1523), .A3(n1522), .A4(n1521), .ZN(n1535) );
  nd04d0 U63 ( .A1(n1842), .A2(n1841), .A3(n1840), .A4(n1839), .ZN(n1853) );
  nd04d0 U64 ( .A1(n1800), .A2(n1799), .A3(n1798), .A4(n1797), .ZN(n1801) );
  nd04d0 U65 ( .A1(n1623), .A2(n1622), .A3(n1621), .A4(n1620), .ZN(n1624) );
  nd04d0 U66 ( .A1(n1145), .A2(n1144), .A3(n1143), .A4(n1142), .ZN(n1157) );
  nd04d0 U67 ( .A1(n1150), .A2(n1149), .A3(n1148), .A4(n1147), .ZN(n1156) );
  nd04d0 U68 ( .A1(n1057), .A2(n1056), .A3(n1055), .A4(n1054), .ZN(n1068) );
  nd04d0 U69 ( .A1(n1083), .A2(n1082), .A3(n1081), .A4(n1080), .ZN(n1089) );
  nd04d0 U70 ( .A1(n1087), .A2(n1086), .A3(n1085), .A4(n1084), .ZN(n1088) );
  nd04d0 U71 ( .A1(n1127), .A2(n1126), .A3(n1125), .A4(n1124), .ZN(n1133) );
  nd04d0 U72 ( .A1(n1061), .A2(n1060), .A3(n1059), .A4(n1058), .ZN(n1067) );
  nd04d0 U73 ( .A1(n1097), .A2(n1096), .A3(n1095), .A4(n1094), .ZN(n1113) );
  nd04d0 U74 ( .A1(n2005), .A2(n2004), .A3(n2003), .A4(n2002), .ZN(n2011) );
  nd04d0 U75 ( .A1(n999), .A2(n998), .A3(n997), .A4(n996), .ZN(n1000) );
  nd04d0 U76 ( .A1(n886), .A2(n885), .A3(n884), .A4(n883), .ZN(n913) );
  nd04d0 U77 ( .A1(n1966), .A2(n1965), .A3(n1964), .A4(n1963), .ZN(n1977) );
  nd04d0 U78 ( .A1(n1243), .A2(n1242), .A3(n1241), .A4(n1240), .ZN(n1244) );
  nd04d0 U79 ( .A1(n1220), .A2(n1219), .A3(n1218), .A4(n1217), .ZN(n1247) );
  nd04d0 U80 ( .A1(n1207), .A2(n1206), .A3(n1205), .A4(n1204), .ZN(n1208) );
  nd04d0 U81 ( .A1(n2026), .A2(n2025), .A3(n2024), .A4(n2023), .ZN(n2027) );
  nd04d0 U82 ( .A1(n991), .A2(n990), .A3(n989), .A4(n988), .ZN(n1002) );
  nd04d0 U83 ( .A1(n1184), .A2(n1183), .A3(n1182), .A4(n1181), .ZN(n1210) );
  nd04d0 U84 ( .A1(n2022), .A2(n2021), .A3(n2020), .A4(n2019), .ZN(n2028) );
  nd04d0 U85 ( .A1(n1230), .A2(n1229), .A3(n1228), .A4(n1227), .ZN(n1245) );
  nd04d0 U86 ( .A1(n1141), .A2(n1140), .A3(n1139), .A4(n1138), .ZN(n1158) );
  nd04d0 U87 ( .A1(n890), .A2(n889), .A3(n888), .A4(n887), .ZN(n912) );
  nd04d0 U88 ( .A1(n896), .A2(n895), .A3(n894), .A4(n893), .ZN(n911) );
  nd04d0 U89 ( .A1(n1065), .A2(n1064), .A3(n1063), .A4(n1062), .ZN(n1066) );
  nd04d0 U90 ( .A1(n2098), .A2(n2097), .A3(n2096), .A4(n2095), .ZN(n2099) );
  nd04d0 U91 ( .A1(n1172), .A2(n1171), .A3(n1170), .A4(n1169), .ZN(n1211) );
  nd04d0 U92 ( .A1(n1109), .A2(n1108), .A3(n1107), .A4(n1106), .ZN(n1110) );
  nd04d0 U93 ( .A1(n1123), .A2(n1122), .A3(n1121), .A4(n1120), .ZN(n1134) );
  nd04d0 U94 ( .A1(n1101), .A2(n1100), .A3(n1099), .A4(n1098), .ZN(n1112) );
  nd04d0 U95 ( .A1(n1131), .A2(n1130), .A3(n1129), .A4(n1128), .ZN(n1132) );
  nd04d0 U96 ( .A1(n1154), .A2(n1153), .A3(n1152), .A4(n1151), .ZN(n1155) );
  nd04d0 U97 ( .A1(n2080), .A2(n2079), .A3(n2078), .A4(n2077), .ZN(n2081) );
  nd04d0 U98 ( .A1(n1599), .A2(n1598), .A3(n1597), .A4(n1596), .ZN(n1626) );
  nd04d0 U99 ( .A1(n1587), .A2(n1586), .A3(n1585), .A4(n1584), .ZN(n1627) );
  nd04d0 U100 ( .A1(n1441), .A2(n1440), .A3(n1439), .A4(n1438), .ZN(n1442) );
  nd04d0 U101 ( .A1(n1404), .A2(n1403), .A3(n1402), .A4(n1401), .ZN(n1415) );
  nd04d0 U102 ( .A1(n1408), .A2(n1407), .A3(n1406), .A4(n1405), .ZN(n1414) );
  nd04d0 U103 ( .A1(n1905), .A2(n1904), .A3(n1903), .A4(n1902), .ZN(n1911) );
  nd04d0 U104 ( .A1(n1528), .A2(n1527), .A3(n1526), .A4(n1525), .ZN(n1534) );
  nd04d0 U105 ( .A1(n1810), .A2(n1809), .A3(n1808), .A4(n1807), .ZN(n1823) );
  nd04d0 U106 ( .A1(n1498), .A2(n1497), .A3(n1496), .A4(n1495), .ZN(n1504) );
  nd04d0 U107 ( .A1(n1558), .A2(n1557), .A3(n1556), .A4(n1555), .ZN(n1565) );
  nd04d0 U108 ( .A1(n1554), .A2(n1553), .A3(n1552), .A4(n1551), .ZN(n1566) );
  nd04d0 U109 ( .A1(n1459), .A2(n1458), .A3(n1457), .A4(n1456), .ZN(n1475) );
  nd04d0 U110 ( .A1(n1827), .A2(n1826), .A3(n1825), .A4(n1824), .ZN(n1838) );
  nd04d0 U111 ( .A1(n1550), .A2(n1549), .A3(n1548), .A4(n1547), .ZN(n1567) );
  nd04d0 U112 ( .A1(n1463), .A2(n1462), .A3(n1461), .A4(n1460), .ZN(n1474) );
  nd04d0 U113 ( .A1(n1318), .A2(n1317), .A3(n1316), .A4(n1315), .ZN(n1329) );
  nd04d0 U114 ( .A1(n1289), .A2(n1288), .A3(n1287), .A4(n1286), .ZN(n1300) );
  nd04d0 U115 ( .A1(n1293), .A2(n1292), .A3(n1291), .A4(n1290), .ZN(n1299) );
  nd04d0 U116 ( .A1(n1985), .A2(n1984), .A3(n1983), .A4(n1982), .ZN(n1991) );
  nd04d0 U117 ( .A1(n1263), .A2(n1262), .A3(n1261), .A4(n1260), .ZN(n1274) );
  nd04d0 U118 ( .A1(n1267), .A2(n1266), .A3(n1265), .A4(n1264), .ZN(n1273) );
  nd04d0 U119 ( .A1(n1224), .A2(n1223), .A3(n1222), .A4(n1221), .ZN(n1246) );
  nd04d0 U120 ( .A1(n1970), .A2(n1969), .A3(n1968), .A4(n1967), .ZN(n1976) );
  nd04d0 U121 ( .A1(n1371), .A2(n1370), .A3(n1369), .A4(n1368), .ZN(n1387) );
  nd04d0 U122 ( .A1(n1888), .A2(n1887), .A3(n1886), .A4(n1885), .ZN(n1889) );
  nd04d0 U123 ( .A1(n1383), .A2(n1382), .A3(n1381), .A4(n1380), .ZN(n1384) );
  nd04d0 U124 ( .A1(n1342), .A2(n1341), .A3(n1340), .A4(n1339), .ZN(n1358) );
  nd04d0 U125 ( .A1(n1346), .A2(n1345), .A3(n1344), .A4(n1343), .ZN(n1357) );
  nd04d0 U126 ( .A1(n1350), .A2(n1349), .A3(n1348), .A4(n1347), .ZN(n1356) );
  nd04d0 U127 ( .A1(n1354), .A2(n1353), .A3(n1352), .A4(n1351), .ZN(n1355) );
  nd04d0 U128 ( .A1(n1862), .A2(n1861), .A3(n1860), .A4(n1859), .ZN(n1874) );
  nd04d0 U129 ( .A1(n2204), .A2(n2203), .A3(n2202), .A4(n2201), .ZN(n2213) );
  nd04d0 U130 ( .A1(n1031), .A2(n1030), .A3(n1029), .A4(n1028), .ZN(n1047) );
  nd04d0 U131 ( .A1(n1039), .A2(n1038), .A3(n1037), .A4(n1036), .ZN(n1045) );
  nd04d0 U132 ( .A1(n2104), .A2(n2103), .A3(n2102), .A4(n2101), .ZN(n2110) );
  nd04d0 U133 ( .A1(n1009), .A2(n1008), .A3(n1007), .A4(n1006), .ZN(n1025) );
  nd04d0 U134 ( .A1(n1013), .A2(n1012), .A3(n1011), .A4(n1010), .ZN(n1024) );
  nd04d0 U135 ( .A1(n1017), .A2(n1016), .A3(n1015), .A4(n1014), .ZN(n1023) );
  nd04d0 U136 ( .A1(n1021), .A2(n1020), .A3(n1019), .A4(n1018), .ZN(n1022) );
  nd04d0 U137 ( .A1(n987), .A2(n986), .A3(n985), .A4(n984), .ZN(n1003) );
  nd04d0 U138 ( .A1(n2118), .A2(n2117), .A3(n2116), .A4(n2115), .ZN(n2128) );
  nd04d0 U139 ( .A1(n995), .A2(n994), .A3(n993), .A4(n992), .ZN(n1001) );
  nd04d0 U140 ( .A1(n965), .A2(n964), .A3(n963), .A4(n962), .ZN(n981) );
  nd04d0 U141 ( .A1(n969), .A2(n968), .A3(n967), .A4(n966), .ZN(n980) );
  nd04d0 U142 ( .A1(n977), .A2(n976), .A3(n975), .A4(n974), .ZN(n978) );
  nd04d0 U143 ( .A1(n951), .A2(n950), .A3(n949), .A4(n948), .ZN(n957) );
  nd04d0 U144 ( .A1(n2229), .A2(n2228), .A3(n2227), .A4(n2226), .ZN(n2250) );
  nd04d0 U145 ( .A1(n1437), .A2(n1436), .A3(n1435), .A4(n1434), .ZN(n1443) );
  nd04d0 U146 ( .A1(n1925), .A2(n1924), .A3(n1923), .A4(n1922), .ZN(n1926) );
  nd04d0 U147 ( .A1(n1831), .A2(n1830), .A3(n1829), .A4(n1828), .ZN(n1837) );
  nd04d0 U148 ( .A1(n1502), .A2(n1501), .A3(n1500), .A4(n1499), .ZN(n1503) );
  nd04d0 U149 ( .A1(n1835), .A2(n1834), .A3(n1833), .A4(n1832), .ZN(n1836) );
  nd04d0 U150 ( .A1(n1490), .A2(n1489), .A3(n1488), .A4(n1487), .ZN(n1506) );
  nd04d0 U151 ( .A1(n1412), .A2(n1411), .A3(n1410), .A4(n1409), .ZN(n1413) );
  nd04d0 U152 ( .A1(n1314), .A2(n1313), .A3(n1312), .A4(n1311), .ZN(n1330) );
  nd04d0 U153 ( .A1(n1611), .A2(n1610), .A3(n1609), .A4(n1608), .ZN(n1625) );
  nd04d0 U154 ( .A1(n2108), .A2(n2107), .A3(n2106), .A4(n2105), .ZN(n2109) );
  nd04d0 U155 ( .A1(n1075), .A2(n1074), .A3(n1073), .A4(n1072), .ZN(n1091) );
  nd04d0 U156 ( .A1(n1105), .A2(n1104), .A3(n1103), .A4(n1102), .ZN(n1111) );
  nd04d0 U157 ( .A1(n947), .A2(n946), .A3(n945), .A4(n944), .ZN(n958) );
  nd04d0 U158 ( .A1(n973), .A2(n972), .A3(n971), .A4(n970), .ZN(n979) );
  nd04d0 U159 ( .A1(n1974), .A2(n1973), .A3(n1972), .A4(n1971), .ZN(n1975) );
  nd04d0 U160 ( .A1(n1297), .A2(n1296), .A3(n1295), .A4(n1294), .ZN(n1298) );
  nd04d0 U161 ( .A1(n1285), .A2(n1284), .A3(n1283), .A4(n1282), .ZN(n1301) );
  nd04d0 U162 ( .A1(n1195), .A2(n1194), .A3(n1193), .A4(n1192), .ZN(n1209) );
  nd04d0 U163 ( .A1(n2009), .A2(n2008), .A3(n2007), .A4(n2006), .ZN(n2010) );
  nd04d0 U164 ( .A1(n1079), .A2(n1078), .A3(n1077), .A4(n1076), .ZN(n1090) );
  nd04d0 U165 ( .A1(n1053), .A2(n1052), .A3(n1051), .A4(n1050), .ZN(n1069) );
  nd04d0 U166 ( .A1(n1043), .A2(n1042), .A3(n1041), .A4(n1040), .ZN(n1044) );
  nd04d0 U167 ( .A1(n1909), .A2(n1908), .A3(n1907), .A4(n1906), .ZN(n1910) );
  nd04d0 U168 ( .A1(n1981), .A2(n1980), .A3(n1979), .A4(n1978), .ZN(n1992) );
  nd03d0 U169 ( .A1(n2044), .A2(n2043), .A3(n2042), .ZN(n2050) );
  nd03d0 U170 ( .A1(n2089), .A2(n2088), .A3(n2087), .ZN(n2090) );
  nd03d0 U171 ( .A1(n2036), .A2(n2035), .A3(n2034), .ZN(n2060) );
  nd03d0 U172 ( .A1(n2018), .A2(n2017), .A3(n2016), .ZN(n2029) );
  nd03d0 U173 ( .A1(n1951), .A2(n1950), .A3(n1949), .ZN(n1952) );
  nd03d0 U174 ( .A1(n1917), .A2(n1916), .A3(n1915), .ZN(n1928) );
  nd03d0 U175 ( .A1(n1794), .A2(n1793), .A3(n1792), .ZN(n1795) );
  nd12d0 U176 ( .A1(n818), .A2(n817), .ZN(n867) );
  or02d0 U177 ( .A1(n831), .A2(n864), .Z(n2262) );
  nd02d0 U178 ( .A1(N865), .A2(n766), .ZN(n699) );
  nd03d0 U179 ( .A1(n784), .A2(n719), .A3(n684), .ZN(n736) );
  nd03d0 U180 ( .A1(N867), .A2(n632), .A3(n631), .ZN(n634) );
  nd02d0 U181 ( .A1(N861), .A2(N860), .ZN(n731) );
  nd03d0 U182 ( .A1(n684), .A2(n665), .A3(N862), .ZN(n786) );
  nd03d0 U183 ( .A1(n1673), .A2(n1696), .A3(n1559), .ZN(n1541) );
  nd03d0 U184 ( .A1(wb_adr_i[25]), .A2(wb_adr_i[29]), .A3(wb_adr_i[26]), .ZN(
        n573) );
  nd03d0 U185 ( .A1(wb_cyc_i), .A2(wb_stb_i), .A3(n566), .ZN(n572) );
  nd12d0 U186 ( .A1(n3169), .A2(n2254), .ZN(n3257) );
  nd03d0 U187 ( .A1(n2137), .A2(n2142), .A3(n1719), .ZN(n827) );
  nd02d0 U188 ( .A1(N864), .A2(n615), .ZN(n778) );
  nd03d0 U189 ( .A1(N862), .A2(n712), .A3(n665), .ZN(n776) );
  nd03d0 U190 ( .A1(N863), .A2(n783), .A3(n707), .ZN(n734) );
  nd02d0 U191 ( .A1(spimemio_flash_io0_oeb), .A2(n2302), .ZN(n3390) );
  inv0d0 U192 ( .I(n3242), .ZN(n475) );
  inv0d1 U193 ( .I(n481), .ZN(n3343) );
  inv0d1 U194 ( .I(n482), .ZN(n3337) );
  inv0d1 U195 ( .I(n482), .ZN(n3379) );
  inv0d1 U196 ( .I(n484), .ZN(n3339) );
  inv0d1 U197 ( .I(n483), .ZN(n3338) );
  inv0d1 U198 ( .I(n484), .ZN(n3336) );
  inv0d1 U199 ( .I(n482), .ZN(n3363) );
  inv0d1 U200 ( .I(n482), .ZN(n3364) );
  inv0d1 U201 ( .I(n482), .ZN(n3365) );
  inv0d1 U202 ( .I(n482), .ZN(n3366) );
  inv0d1 U203 ( .I(n483), .ZN(n3371) );
  inv0d1 U204 ( .I(n483), .ZN(n3368) );
  inv0d1 U205 ( .I(n483), .ZN(n3369) );
  inv0d1 U206 ( .I(n483), .ZN(n3370) );
  inv0d1 U207 ( .I(n482), .ZN(n3355) );
  inv0d1 U208 ( .I(n481), .ZN(n3356) );
  inv0d1 U209 ( .I(n484), .ZN(n3357) );
  inv0d1 U210 ( .I(n483), .ZN(n3358) );
  inv0d1 U211 ( .I(n482), .ZN(n3348) );
  inv0d1 U212 ( .I(n483), .ZN(n3349) );
  inv0d1 U213 ( .I(n482), .ZN(n3350) );
  inv0d1 U214 ( .I(n483), .ZN(n3351) );
  inv0d1 U215 ( .I(n482), .ZN(n3377) );
  inv0d1 U216 ( .I(n483), .ZN(n3382) );
  inv0d1 U217 ( .I(n482), .ZN(n3386) );
  inv0d1 U218 ( .I(n483), .ZN(n3381) );
  inv0d1 U219 ( .I(n484), .ZN(n3378) );
  inv0d1 U220 ( .I(n484), .ZN(n3383) );
  inv0d1 U221 ( .I(n484), .ZN(n3387) );
  inv0d1 U222 ( .I(n484), .ZN(n3375) );
  inv0d1 U223 ( .I(n481), .ZN(n3380) );
  inv0d1 U224 ( .I(n481), .ZN(n3384) );
  inv0d1 U225 ( .I(n481), .ZN(n3385) );
  inv0d1 U226 ( .I(n481), .ZN(n3376) );
  inv0d1 U227 ( .I(n483), .ZN(n3345) );
  inv0d1 U228 ( .I(n481), .ZN(n3346) );
  inv0d1 U229 ( .I(n481), .ZN(n3347) );
  inv0d1 U230 ( .I(n3257), .ZN(n3258) );
  inv0d2 U231 ( .I(wbbd_busy), .ZN(n2341) );
  nr02d2 U232 ( .A1(n862), .A2(n825), .ZN(n2264) );
  buffd3 U233 ( .I(n1785), .Z(n1778) );
  inv0d1 U234 ( .I(n1214), .ZN(n1632) );
  inv0d1 U235 ( .I(n2262), .ZN(n2094) );
  aoim22d1 U236 ( .A1(n828), .A2(n863), .B1(serial_bb_data_1), .B2(n828), .Z(
        n3038) );
  inv0d1 U237 ( .I(n827), .ZN(n828) );
  inv0d1 U238 ( .I(n822), .ZN(n824) );
  inv0d2 U239 ( .I(n3237), .ZN(n863) );
  nr02d2 U240 ( .A1(n843), .A2(n867), .ZN(n844) );
  inv0d2 U241 ( .I(n3236), .ZN(n1782) );
  inv0d2 U242 ( .I(n2333), .ZN(n3228) );
  inv0d2 U243 ( .I(n3235), .ZN(n1786) );
  inv0d2 U244 ( .I(wb_rstn_i), .ZN(n3292) );
  inv0d1 U245 ( .I(n482), .ZN(n3340) );
  inv0d2 U246 ( .I(n1649), .ZN(serial_clock) );
  nd02d0 U247 ( .A1(spi_is_enabled), .A2(n497), .ZN(n2342) );
  nd04d0 U248 ( .A1(n2048), .A2(n2047), .A3(n2046), .A4(n2045), .ZN(n2049) );
  nd03d0 U249 ( .A1(n2032), .A2(n2031), .A3(n2030), .ZN(n2033) );
  nd04d0 U250 ( .A1(n2125), .A2(n2124), .A3(n2123), .A4(n2122), .ZN(n2126) );
  nd03d0 U251 ( .A1(n2121), .A2(n2120), .A3(n2119), .ZN(n2127) );
  nd04d0 U252 ( .A1(n1989), .A2(n1988), .A3(n1987), .A4(n1986), .ZN(n1990) );
  nd03d0 U253 ( .A1(n1682), .A2(n1676), .A3(n1672), .ZN(n1225) );
  nd03d0 U254 ( .A1(n1679), .A2(n1673), .A3(n1683), .ZN(n1231) );
  nd04d0 U255 ( .A1(n2210), .A2(n2209), .A3(n2208), .A4(n2207), .ZN(n2212) );
  nd04d0 U256 ( .A1(n2154), .A2(n2153), .A3(n2152), .A4(n2151), .ZN(n2155) );
  nd04d0 U257 ( .A1(n2040), .A2(n2039), .A3(n2038), .A4(n2037), .ZN(n2059) );
  nd04d0 U258 ( .A1(n1921), .A2(n1920), .A3(n1919), .A4(n1918), .ZN(n1927) );
  nd04d0 U259 ( .A1(n1846), .A2(n1845), .A3(n1844), .A4(n1843), .ZN(n1852) );
  nr02d0 U260 ( .A1(N864), .A2(N865), .ZN(n632) );
  nr02d0 U261 ( .A1(n741), .A2(n629), .ZN(n722) );
  nd04d0 U262 ( .A1(n2246), .A2(n2245), .A3(n2244), .A4(n2243), .ZN(n2248) );
  nr03d0 U263 ( .A1(n2029), .A2(n2028), .A3(n2027), .ZN(n2063) );
  nr04d0 U264 ( .A1(n1953), .A2(n1928), .A3(n1927), .A4(n1926), .ZN(n1929) );
  nr04d0 U265 ( .A1(wb_adr_i[24]), .A2(wb_adr_i[16]), .A3(wb_adr_i[13]), .A4(
        wb_adr_i[15]), .ZN(n567) );
  nr04d0 U266 ( .A1(n748), .A2(n769), .A3(n747), .A4(n746), .ZN(n749) );
  nd04d0 U267 ( .A1(n2194), .A2(n2193), .A3(n2192), .A4(n2191), .ZN(n2219) );
  nd04d0 U268 ( .A1(n1806), .A2(n1805), .A3(n1804), .A4(n1803), .ZN(n1858) );
  nd04d0 U269 ( .A1(n1532), .A2(n1531), .A3(n1530), .A4(n1529), .ZN(n1533) );
  nd04d0 U270 ( .A1(n1467), .A2(n1466), .A3(n1465), .A4(n1464), .ZN(n1473) );
  nd04d0 U271 ( .A1(n1400), .A2(n1399), .A3(n1398), .A4(n1397), .ZN(n1416) );
  nd04d0 U272 ( .A1(n1326), .A2(n1325), .A3(n1324), .A4(n1323), .ZN(n1327) );
  nd04d0 U273 ( .A1(n1271), .A2(n1270), .A3(n1269), .A4(n1268), .ZN(n1272) );
  nd04d0 U274 ( .A1(n909), .A2(n908), .A3(n907), .A4(n906), .ZN(n910) );
  nd04d0 U275 ( .A1(n1119), .A2(n1118), .A3(n1117), .A4(n1116), .ZN(n1135) );
  nd04d0 U276 ( .A1(n1035), .A2(n1034), .A3(n1033), .A4(n1032), .ZN(n1046) );
  nd04d0 U277 ( .A1(n955), .A2(n954), .A3(n953), .A4(n952), .ZN(n956) );
  nr02d0 U278 ( .A1(n741), .A2(n699), .ZN(n712) );
  nd04d0 U279 ( .A1(n677), .A2(n676), .A3(n690), .A4(n675), .ZN(n678) );
  nr02d0 U280 ( .A1(n630), .A2(n744), .ZN(n680) );
  nr02d0 U281 ( .A1(n552), .A2(n551), .ZN(n556) );
  nd12d0 U282 ( .A1(n839), .A2(n2255), .ZN(n3206) );
  nd12d0 U283 ( .A1(n3169), .A2(n2276), .ZN(n3118) );
  nr02d0 U284 ( .A1(n1740), .A2(n1758), .ZN(n1739) );
  nr02d0 U285 ( .A1(n633), .A2(n1758), .ZN(n1717) );
  nr04d0 U286 ( .A1(n1475), .A2(n1474), .A3(n1473), .A4(n1472), .ZN(n1486) );
  nr04d0 U287 ( .A1(n1301), .A2(n1300), .A3(n1299), .A4(n1298), .ZN(n1310) );
  nr04d0 U288 ( .A1(n1113), .A2(n1112), .A3(n1111), .A4(n1110), .ZN(n1115) );
  nr04d0 U289 ( .A1(n959), .A2(n958), .A3(n957), .A4(n956), .ZN(n961) );
  nr04d0 U290 ( .A1(wb_adr_i[30]), .A2(n573), .A3(n572), .A4(n571), .ZN(n812)
         );
  nr02d0 U291 ( .A1(n1896), .A2(n872), .ZN(n3209) );
  nr02d0 U292 ( .A1(n1815), .A2(n872), .ZN(n3192) );
  nr02d0 U293 ( .A1(n2072), .A2(n1711), .ZN(n3143) );
  nr02d0 U294 ( .A1(irq[0]), .A2(n1706), .ZN(n1704) );
  nr02d0 U295 ( .A1(n2262), .A2(n872), .ZN(n3105) );
  nd12d0 U296 ( .A1(n563), .A2(n555), .ZN(n512) );
  nd12d0 U297 ( .A1(n806), .A2(n487), .ZN(n3058) );
  nr02d0 U298 ( .A1(wbbd_sck), .A2(n2341), .ZN(n2340) );
  inv0d0 U299 ( .I(\hkspi/addr[1] ), .ZN(n526) );
  inv0d0 U300 ( .I(\hkspi/state[1] ), .ZN(n517) );
  inv0d0 U301 ( .I(\hkspi/state[2] ), .ZN(n500) );
  nd03d0 U302 ( .A1(\hkspi/state[0] ), .A2(n517), .A3(n500), .ZN(n523) );
  nd02d0 U303 ( .A1(n2341), .A2(n523), .ZN(n485) );
  inv0d0 U304 ( .I(wbbd_addr[1]), .ZN(n657) );
  inv0d0 U305 ( .I(\hkspi/addr[0] ), .ZN(n527) );
  inv0d1 U306 ( .I(n523), .ZN(n555) );
  nd02d0 U307 ( .A1(n2341), .A2(n555), .ZN(n486) );
  oai222d1 U308 ( .A1(n526), .A2(n485), .B1(n657), .B2(n2341), .C1(n527), .C2(
        n486), .ZN(n817) );
  inv0d0 U309 ( .I(\hkspi/addr[2] ), .ZN(n529) );
  inv0d0 U310 ( .I(wbbd_addr[2]), .ZN(n692) );
  oai222d1 U311 ( .A1(n529), .A2(n485), .B1(n692), .B2(n2341), .C1(n526), .C2(
        n486), .ZN(n818) );
  nd12d0 U312 ( .A1(n817), .A2(n818), .ZN(n864) );
  inv0d0 U313 ( .I(\hkspi/addr[3] ), .ZN(n535) );
  aoi22d1 U314 ( .A1(n555), .A2(n529), .B1(n535), .B2(n523), .ZN(n476) );
  aoi22d1 U315 ( .A1(wbbd_busy), .A2(wbbd_addr[3]), .B1(n476), .B2(n2341), 
        .ZN(n829) );
  inv0d0 U316 ( .I(n829), .ZN(n816) );
  aoi22d1 U317 ( .A1(n555), .A2(\hkspi/addr[5] ), .B1(\hkspi/addr[6] ), .B2(
        n523), .ZN(n477) );
  aoim22d1 U318 ( .A1(n477), .A2(n2341), .B1(n2341), .B2(wbbd_addr[6]), .Z(
        n830) );
  nd02d0 U319 ( .A1(n816), .A2(n830), .ZN(n832) );
  aoim22d1 U320 ( .A1(n555), .A2(n535), .B1(\hkspi/addr[4] ), .B2(n555), .Z(
        n478) );
  aoi22d1 U321 ( .A1(wbbd_busy), .A2(wbbd_addr[4]), .B1(n478), .B2(n2341), 
        .ZN(n861) );
  nd12d0 U322 ( .A1(n832), .A2(n861), .ZN(n825) );
  nr02d0 U323 ( .A1(n864), .A2(n825), .ZN(n2268) );
  buffd1 U324 ( .I(n2268), .Z(n2195) );
  inv0d0 U325 ( .I(n486), .ZN(n480) );
  inv0d0 U326 ( .I(n485), .ZN(n479) );
  aoi222d1 U327 ( .A1(wbbd_busy), .A2(wbbd_addr[0]), .B1(n480), .B2(idata[0]), 
        .C1(n479), .C2(\hkspi/addr[0] ), .ZN(n813) );
  inv0d0 U328 ( .I(n813), .ZN(n814) );
  aoi222d1 U329 ( .A1(wbbd_busy), .A2(wbbd_addr[5]), .B1(n480), .B2(
        \hkspi/addr[4] ), .C1(n479), .C2(\hkspi/addr[5] ), .ZN(n815) );
  nr02d0 U330 ( .A1(n814), .A2(n815), .ZN(n2211) );
  nd02d0 U331 ( .A1(n2195), .A2(n2211), .ZN(n1740) );
  inv0d0 U332 ( .I(n1740), .ZN(n620) );
  nr02d0 U333 ( .A1(pass_thru_mgmt_delay), .A2(n3387), .ZN(pad_flash_csb_oeb)
         );
  nr02d0 U334 ( .A1(pass_thru_mgmt), .A2(n3383), .ZN(pad_flash_clk_oeb) );
  inv0d0 U335 ( .I(mgmt_gpio_in[4]), .ZN(n3296) );
  buffd1 U336 ( .I(csclk), .Z(n3322) );
  buffd1 U337 ( .I(n3322), .Z(n3303) );
  buffd1 U338 ( .I(n3303), .Z(n3329) );
  buffd1 U339 ( .I(n3329), .Z(n3319) );
  buffd1 U340 ( .I(n3319), .Z(n3323) );
  buffd1 U341 ( .I(n3323), .Z(n3326) );
  buffd1 U342 ( .I(n3326), .Z(n3311) );
  buffd1 U343 ( .I(n3323), .Z(n3305) );
  buffd1 U344 ( .I(n3305), .Z(n3328) );
  buffd1 U345 ( .I(n3328), .Z(n3318) );
  buffd1 U346 ( .I(n3323), .Z(n3327) );
  buffd1 U347 ( .I(n3327), .Z(n3308) );
  buffd1 U348 ( .I(mgmt_gpio_in[4]), .Z(n3291) );
  buffd1 U349 ( .I(n3323), .Z(n3307) );
  buffd1 U350 ( .I(n3307), .Z(n3325) );
  buffd1 U351 ( .I(n3325), .Z(n3310) );
  buffd1 U352 ( .I(n3325), .Z(n3309) );
  buffd1 U353 ( .I(wb_clk_i), .Z(n3331) );
  buffd1 U354 ( .I(wb_clk_i), .Z(n3332) );
  buffd1 U355 ( .I(wb_clk_i), .Z(n3330) );
  buffd1 U356 ( .I(wb_clk_i), .Z(n3333) );
  buffd1 U357 ( .I(n3323), .Z(n3298) );
  buffd1 U358 ( .I(n3323), .Z(n3314) );
  buffd1 U359 ( .I(n3314), .Z(n3321) );
  buffd1 U360 ( .I(n3321), .Z(n3324) );
  buffd1 U361 ( .I(n3324), .Z(n3300) );
  buffd1 U362 ( .I(n3322), .Z(n3304) );
  buffd1 U363 ( .I(n3307), .Z(n3302) );
  buffd1 U364 ( .I(n3321), .Z(n3297) );
  buffd1 U365 ( .I(n3297), .Z(n3301) );
  buffd1 U366 ( .I(n3303), .Z(n3320) );
  buffd3 U367 ( .I(n3320), .Z(n3312) );
  buffd1 U368 ( .I(n3312), .Z(n3316) );
  buffd1 U369 ( .I(n3303), .Z(n3313) );
  buffd1 U370 ( .I(n3323), .Z(n3306) );
  buffd1 U371 ( .I(n3306), .Z(n3315) );
  buffd1 U372 ( .I(n3306), .Z(n3317) );
  buffd1 U373 ( .I(n3323), .Z(n3299) );
  buffd1 U374 ( .I(wb_clk_i), .Z(n3334) );
  inv0d0 U375 ( .I(porb), .ZN(n481) );
  buffd1 U376 ( .I(n481), .Z(n482) );
  inv0d0 U377 ( .I(n482), .ZN(n3367) );
  buffd1 U378 ( .I(n481), .Z(n483) );
  inv0d0 U379 ( .I(n482), .ZN(n3359) );
  inv0d0 U380 ( .I(n483), .ZN(n3360) );
  inv0d0 U381 ( .I(n482), .ZN(n3361) );
  inv0d0 U382 ( .I(n482), .ZN(n3362) );
  inv0d0 U383 ( .I(n483), .ZN(n3372) );
  inv0d0 U384 ( .I(n483), .ZN(n3373) );
  inv0d0 U385 ( .I(n483), .ZN(n3374) );
  inv0d0 U386 ( .I(porb), .ZN(n484) );
  nr02d1 U387 ( .A1(\_1_net_[0] ), .A2(n484), .ZN(n2523) );
  buffd1 U388 ( .I(n2523), .Z(n3294) );
  buffd1 U389 ( .I(n2523), .Z(n3295) );
  buffd1 U390 ( .I(n2523), .Z(n3293) );
  inv0d0 U391 ( .I(n483), .ZN(n3341) );
  inv0d0 U392 ( .I(n484), .ZN(n3342) );
  inv0d0 U393 ( .I(n483), .ZN(n3344) );
  inv0d0 U394 ( .I(n482), .ZN(n3352) );
  inv0d0 U395 ( .I(n483), .ZN(n3353) );
  inv0d0 U396 ( .I(n484), .ZN(n3354) );
  inv0d0 U397 ( .I(serial_bb_enable), .ZN(n2181) );
  mx02d1 U398 ( .I0(serial_bb_resetn), .I1(serial_resetn_pre), .S(n2181), .Z(
        serial_resetn) );
  nr02d0 U399 ( .A1(n829), .A2(n830), .ZN(n853) );
  inv0d0 U400 ( .I(n861), .ZN(n834) );
  nd02d0 U401 ( .A1(n853), .A2(n834), .ZN(n843) );
  or02d0 U402 ( .A1(n818), .A2(n817), .Z(n871) );
  nr02d1 U403 ( .A1(n843), .A2(n871), .ZN(n2236) );
  inv0d0 U404 ( .I(n2236), .ZN(n1898) );
  aoi22d1 U405 ( .A1(wbbd_busy), .A2(wbbd_write), .B1(wrstb), .B2(n2341), .ZN(
        n1705) );
  inv0d0 U406 ( .I(\hkspi/addr[6] ), .ZN(n554) );
  inv0d0 U407 ( .I(\hkspi/addr[7] ), .ZN(n558) );
  oai22d1 U408 ( .A1(n554), .A2(n486), .B1(n485), .B2(n558), .ZN(n819) );
  nr02d0 U409 ( .A1(n1705), .A2(n819), .ZN(n1719) );
  nd02d1 U410 ( .A1(n2211), .A2(n1719), .ZN(n874) );
  nr02d1 U411 ( .A1(n1898), .A2(n874), .ZN(n3164) );
  aoi22d1 U412 ( .A1(wbbd_busy), .A2(wbbd_data[2]), .B1(idata[2]), .B2(n2341), 
        .ZN(n849) );
  aoim22d1 U413 ( .A1(n3164), .A2(n849), .B1(\gpio_configure[13][2] ), .B2(
        n3164), .Z(n2787) );
  nr02d0 U414 ( .A1(n843), .A2(n864), .ZN(n2068) );
  buffd1 U415 ( .I(n2068), .Z(n2223) );
  inv0d0 U416 ( .I(n2223), .ZN(n1877) );
  nr02d1 U417 ( .A1(n1877), .A2(n874), .ZN(n2326) );
  aoim22d1 U418 ( .A1(n2326), .A2(n849), .B1(\gpio_configure[15][2] ), .B2(
        n2326), .Z(n2807) );
  inv0d0 U419 ( .I(\gpio_configure[36][3] ), .ZN(mgmt_gpio_oeb[36]) );
  inv0d0 U420 ( .I(n2195), .ZN(n2093) );
  nr02d0 U421 ( .A1(n813), .A2(n815), .ZN(n2131) );
  inv0d0 U422 ( .I(n2131), .ZN(n2054) );
  nr02d0 U423 ( .A1(n2093), .A2(n2054), .ZN(n2284) );
  inv0d0 U424 ( .I(n2284), .ZN(n633) );
  inv0d0 U425 ( .I(mgmt_gpio_data_9), .ZN(n2319) );
  nr02d0 U426 ( .A1(\gpio_configure[3][3] ), .A2(hkspi_disable), .ZN(
        spi_is_enabled) );
  inv0d0 U427 ( .I(mgmt_gpio_in[3]), .ZN(n497) );
  inv0d0 U428 ( .I(pass_thru_user), .ZN(n2335) );
  an02d0 U429 ( .A1(mgmt_gpio_in[0]), .A2(debug_mode), .Z(debug_in) );
  inv0d0 U430 ( .I(wbbd_state[3]), .ZN(n581) );
  nr03d0 U431 ( .A1(wbbd_state[2]), .A2(wbbd_state[0]), .A3(n581), .ZN(n806)
         );
  nd02d1 U432 ( .A1(n581), .A2(wbbd_state[0]), .ZN(n797) );
  inv0d0 U433 ( .I(wbbd_state[2]), .ZN(n3277) );
  inv0d0 U434 ( .I(wbbd_state[1]), .ZN(n579) );
  nd02d0 U435 ( .A1(n3277), .A2(n579), .ZN(n803) );
  oai211d1 U436 ( .C1(wbbd_sck), .C2(n581), .A(n797), .B(n803), .ZN(n487) );
  inv0d0 U437 ( .I(pad_flash_io1_di), .ZN(n496) );
  nr02d0 U438 ( .A1(pass_thru_mgmt), .A2(n496), .ZN(spimemio_flash_io1_di) );
  inv0d0 U439 ( .I(\gpio_configure[37][3] ), .ZN(mgmt_gpio_oeb[37]) );
  inv0d0 U440 ( .I(pass_thru_mgmt_delay), .ZN(n2302) );
  mx02d1 U441 ( .I0(idata[0]), .I1(spimemio_flash_io0_do), .S(n2302), .Z(
        pad_flash_io0_do) );
  inv0d0 U442 ( .I(n3390), .ZN(pad_flash_io0_oeb) );
  inv0d0 U443 ( .I(mgmt_gpio_data_13), .ZN(n1751) );
  nr02d0 U444 ( .A1(trap_output_dest), .A2(n1751), .ZN(mgmt_gpio_out[13]) );
  or03d0 U445 ( .A1(reset_reg), .A2(pass_thru_mgmt_delay), .A3(
        \hkspi/pre_pass_thru_mgmt ), .Z(reset) );
  mx02d1 U446 ( .I0(mgmt_gpio_data_15), .I1(user_clock), .S(clk2_output_dest), 
        .Z(mgmt_gpio_out_15_prebuff) );
  inv0d0 U447 ( .I(\gpio_configure[0][3] ), .ZN(n879) );
  mx02d1 U448 ( .I0(n879), .I1(debug_oeb), .S(debug_mode), .Z(mgmt_gpio_oeb[0]) );
  aoim22d1 U449 ( .A1(clk1_output_dest), .A2(n2322), .B1(mgmt_gpio_data_14), 
        .B2(clk1_output_dest), .Z(mgmt_gpio_out_14_prebuff) );
  inv0d0 U450 ( .I(spi_enabled), .ZN(n499) );
  mx02d1 U451 ( .I0(spi_sck), .I1(mgmt_gpio_data_32), .S(n499), .Z(
        mgmt_gpio_out[32]) );
  mx02d1 U452 ( .I0(mgmt_gpio_data_6), .I1(ser_tx), .S(uart_enabled), .Z(
        mgmt_gpio_out[6]) );
  mx02d1 U453 ( .I0(spi_sdo), .I1(mgmt_gpio_data[35]), .S(n499), .Z(
        mgmt_gpio_out[35]) );
  inv0d0 U454 ( .I(idata[0]), .ZN(n2307) );
  inv0d0 U455 ( .I(mgmt_gpio_data_10), .ZN(n1744) );
  inv0d0 U456 ( .I(pass_thru_user_delay), .ZN(n2304) );
  aoi22d1 U457 ( .A1(pass_thru_user_delay), .A2(n2307), .B1(n1744), .B2(n2304), 
        .ZN(mgmt_gpio_out[10]) );
  an02d0 U458 ( .A1(irq_1_inputsrc), .A2(mgmt_gpio_in[7]), .Z(irq[1]) );
  an02d0 U459 ( .A1(irq_2_inputsrc), .A2(mgmt_gpio_in[12]), .Z(irq[2]) );
  nr02d0 U460 ( .A1(\hkspi/state[2] ), .A2(\hkspi/state[0] ), .ZN(n488) );
  nd02d0 U461 ( .A1(\hkspi/state[1] ), .A2(n488), .ZN(n2312) );
  nd03d0 U462 ( .A1(\hkspi/count[2] ), .A2(\hkspi/count[1] ), .A3(
        \hkspi/count[0] ), .ZN(n563) );
  nr02d0 U463 ( .A1(n2312), .A2(n563), .ZN(n521) );
  inv0d0 U464 ( .I(\hkspi/fixed[1] ), .ZN(n515) );
  inv0d0 U465 ( .I(\hkspi/fixed[0] ), .ZN(n511) );
  nd04d0 U466 ( .A1(\hkspi/fixed[2] ), .A2(n521), .A3(n515), .A4(n511), .ZN(
        n513) );
  inv0d0 U467 ( .I(\hkspi/count[2] ), .ZN(n504) );
  inv0d0 U468 ( .I(\hkspi/count[1] ), .ZN(n507) );
  nd02d0 U469 ( .A1(n488), .A2(n517), .ZN(n2316) );
  inv0d0 U470 ( .I(\hkspi/count[0] ), .ZN(n2317) );
  aoi21d1 U471 ( .B1(n2317), .B2(n507), .A(n504), .ZN(n489) );
  aoi211d1 U472 ( .C1(n504), .C2(n507), .A(n2316), .B(n489), .ZN(n516) );
  oan211d1 U473 ( .C1(\hkspi/fixed[2] ), .C2(\hkspi/fixed[1] ), .B(n521), .A(
        n516), .ZN(n491) );
  oai22d1 U474 ( .A1(\hkspi/fixed[1] ), .A2(n516), .B1(\hkspi/fixed[0] ), .B2(
        n491), .ZN(n490) );
  nd02d0 U475 ( .A1(n513), .A2(n490), .ZN(n3094) );
  aoi22d1 U476 ( .A1(idata[0]), .A2(n516), .B1(\hkspi/fixed[0] ), .B2(n491), 
        .ZN(n493) );
  oai211d1 U477 ( .C1(\hkspi/fixed[2] ), .C2(\hkspi/fixed[1] ), .A(n521), .B(
        n511), .ZN(n492) );
  nd02d0 U478 ( .A1(n493), .A2(n492), .ZN(n3095) );
  an02d0 U479 ( .A1(mgmt_gpio_in[5]), .A2(uart_enabled), .Z(ser_rx) );
  an02d0 U480 ( .A1(mgmt_gpio_in[34]), .A2(spi_enabled), .Z(spi_sdi) );
  oai22d1 U481 ( .A1(n2181), .A2(serial_bb_clock), .B1(serial_clock_pre), .B2(
        serial_bb_enable), .ZN(n1649) );
  inv0d0 U482 ( .I(wb_rstn_i), .ZN(n3388) );
  inv0d0 U483 ( .I(n2342), .ZN(n1718) );
  inv0d0 U484 ( .I(sdo), .ZN(n2297) );
  inv0d0 U485 ( .I(mgmt_gpio_data_1), .ZN(n1722) );
  aoi22d1 U486 ( .A1(n1718), .A2(n2297), .B1(n1722), .B2(n2342), .ZN(n494) );
  aoi22d1 U487 ( .A1(pass_thru_user), .A2(mgmt_gpio_in[11]), .B1(n494), .B2(
        n2335), .ZN(n495) );
  inv0d0 U488 ( .I(pass_thru_mgmt), .ZN(n518) );
  aoi22d1 U489 ( .A1(pass_thru_mgmt), .A2(n496), .B1(n495), .B2(n518), .ZN(
        mgmt_gpio_out[1]) );
  inv0d0 U490 ( .I(mgmt_gpio_data_8), .ZN(n1742) );
  aoi22d1 U491 ( .A1(pass_thru_user_delay), .A2(n497), .B1(n1742), .B2(n2304), 
        .ZN(mgmt_gpio_out[8]) );
  inv0d0 U492 ( .I(mgmt_gpio_data_33), .ZN(n823) );
  nd02d0 U493 ( .A1(spi_enabled), .A2(spi_csb), .ZN(n498) );
  oai21d1 U494 ( .B1(spi_enabled), .B2(n823), .A(n498), .ZN(mgmt_gpio_out[33])
         );
  aoi22d1 U495 ( .A1(spi_enabled), .A2(spi_csb), .B1(\gpio_configure[35][3] ), 
        .B2(n499), .ZN(mgmt_gpio_oeb[35]) );
  inv0d0 U496 ( .I(mgmt_gpio_data_0), .ZN(n1721) );
  nr02d0 U497 ( .A1(debug_mode), .A2(n1721), .ZN(mgmt_gpio_out[0]) );
  inv0d0 U498 ( .I(n2312), .ZN(n2315) );
  nd02d0 U499 ( .A1(\hkspi/readmode ), .A2(n2315), .ZN(n2178) );
  inv0d0 U500 ( .I(n2178), .ZN(n2296) );
  aoi21d1 U501 ( .B1(\hkspi/state[2] ), .B2(n517), .A(n2296), .ZN(\hkspi/N34 )
         );
  inv0d0 U502 ( .I(\gpio_configure[1][3] ), .ZN(n877) );
  mx02d1 U503 ( .I0(sdo_enb), .I1(n877), .S(n2342), .Z(mgmt_gpio_oeb[1]) );
  inv0d0 U504 ( .I(\hkspi/pre_pass_thru_mgmt ), .ZN(n509) );
  inv0d0 U505 ( .I(\hkspi/pre_pass_thru_user ), .ZN(n501) );
  nr02d0 U506 ( .A1(n504), .A2(n2316), .ZN(n510) );
  nd03d0 U507 ( .A1(\hkspi/count[1] ), .A2(\hkspi/count[0] ), .A3(n510), .ZN(
        n2303) );
  aon211d1 U508 ( .C1(n509), .C2(n501), .B(n2303), .A(n500), .ZN(n3103) );
  aoi21d1 U509 ( .B1(\hkspi/state[1] ), .B2(\hkspi/state[0] ), .A(
        \hkspi/state[2] ), .ZN(n562) );
  nd02d0 U510 ( .A1(\hkspi/count[0] ), .A2(n562), .ZN(n506) );
  nd03d0 U511 ( .A1(\hkspi/count[1] ), .A2(n510), .A3(n506), .ZN(n2301) );
  nd03d0 U512 ( .A1(\hkspi/count[1] ), .A2(n510), .A3(n509), .ZN(n2300) );
  nd03d0 U513 ( .A1(n2301), .A2(\hkspi/pre_pass_thru_user ), .A3(n2300), .ZN(
        n502) );
  oai21d1 U514 ( .B1(n2301), .B2(n2307), .A(n502), .ZN(n3102) );
  oai21d1 U515 ( .B1(n523), .B2(n563), .A(\hkspi/state[0] ), .ZN(n503) );
  aon211d1 U516 ( .C1(\hkspi/pre_pass_thru_user ), .C2(n509), .B(n2303), .A(
        n503), .ZN(n3101) );
  inv0d0 U517 ( .I(n506), .ZN(n2299) );
  aoim21d1 U518 ( .B1(n562), .B2(\hkspi/count[0] ), .A(n2299), .ZN(n3100) );
  nr02d0 U520 ( .A1(n507), .A2(n506), .ZN(n505) );
  mx02d1 U521 ( .I0(\hkspi/count[2] ), .I1(n504), .S(n505), .Z(n3099) );
  aoi21d1 U522 ( .B1(n507), .B2(n506), .A(n505), .ZN(n3098) );
  nd04d0 U523 ( .A1(idata[0]), .A2(\hkspi/count[0] ), .A3(n510), .A4(n507), 
        .ZN(n508) );
  aon211d1 U524 ( .C1(\hkspi/count[0] ), .C2(n510), .B(n509), .A(n508), .ZN(
        n3097) );
  nr03d0 U525 ( .A1(\hkspi/fixed[2] ), .A2(\hkspi/fixed[1] ), .A3(n511), .ZN(
        n522) );
  aon211d1 U526 ( .C1(n521), .C2(n522), .B(n517), .A(n512), .ZN(n3096) );
  oai21d1 U527 ( .B1(\hkspi/fixed[2] ), .B2(n516), .A(n513), .ZN(n514) );
  aoi21d1 U528 ( .B1(n516), .B2(n515), .A(n514), .ZN(n3093) );
  nd02d0 U529 ( .A1(\hkspi/state[2] ), .A2(n517), .ZN(n519) );
  oai21d1 U530 ( .B1(\hkspi/state[0] ), .B2(n519), .A(n2335), .ZN(n3092) );
  inv0d0 U531 ( .I(\hkspi/state[0] ), .ZN(n520) );
  oai21d1 U532 ( .B1(n520), .B2(n519), .A(n518), .ZN(n3091) );
  inv0d0 U533 ( .I(n521), .ZN(n564) );
  nr02d0 U534 ( .A1(n522), .A2(n564), .ZN(n538) );
  inv0d0 U535 ( .I(n538), .ZN(n552) );
  nd02d0 U536 ( .A1(n523), .A2(n552), .ZN(n547) );
  inv0d0 U537 ( .I(n547), .ZN(n549) );
  aoi21d1 U538 ( .B1(n538), .B2(n527), .A(n549), .ZN(n531) );
  nd02d0 U539 ( .A1(n538), .A2(n526), .ZN(n530) );
  oaim21d1 U540 ( .B1(n523), .B2(n530), .A(\hkspi/addr[0] ), .ZN(n524) );
  oai21d1 U541 ( .B1(n531), .B2(n526), .A(n524), .ZN(n3090) );
  aoi22d1 U542 ( .A1(n555), .A2(idata[0]), .B1(\hkspi/addr[0] ), .B2(n549), 
        .ZN(n525) );
  oai21d1 U543 ( .B1(\hkspi/addr[0] ), .B2(n552), .A(n525), .ZN(n3089) );
  nr03d0 U544 ( .A1(n527), .A2(n529), .A3(n526), .ZN(n533) );
  nr02d0 U545 ( .A1(n533), .A2(n552), .ZN(n532) );
  aon211d1 U546 ( .C1(\hkspi/addr[0] ), .C2(n532), .B(n555), .A(
        \hkspi/addr[1] ), .ZN(n528) );
  aon211d1 U547 ( .C1(n531), .C2(n530), .B(n529), .A(n528), .ZN(n3088) );
  inv0d0 U548 ( .I(n532), .ZN(n536) );
  nd02d0 U549 ( .A1(\hkspi/addr[3] ), .A2(n533), .ZN(n542) );
  inv0d0 U550 ( .I(n542), .ZN(n537) );
  nr02d0 U551 ( .A1(n537), .A2(n552), .ZN(n539) );
  aoi22d1 U552 ( .A1(n555), .A2(\hkspi/addr[2] ), .B1(n533), .B2(n539), .ZN(
        n534) );
  aon211d1 U553 ( .C1(n547), .C2(n536), .B(n535), .A(n534), .ZN(n3087) );
  nd02d0 U554 ( .A1(\hkspi/addr[4] ), .A2(n537), .ZN(n543) );
  nd02d0 U555 ( .A1(n538), .A2(n543), .ZN(n546) );
  nd02d0 U556 ( .A1(n555), .A2(\hkspi/addr[3] ), .ZN(n541) );
  oai21d1 U557 ( .B1(n549), .B2(n539), .A(\hkspi/addr[4] ), .ZN(n540) );
  oai211d1 U558 ( .C1(n542), .C2(n546), .A(n541), .B(n540), .ZN(n3086) );
  inv0d0 U559 ( .I(\hkspi/addr[5] ), .ZN(n545) );
  inv0d0 U560 ( .I(n543), .ZN(n550) );
  aoi21d1 U561 ( .B1(\hkspi/addr[5] ), .B2(n550), .A(n552), .ZN(n548) );
  aoi22d1 U562 ( .A1(n555), .A2(\hkspi/addr[4] ), .B1(n550), .B2(n548), .ZN(
        n544) );
  aon211d1 U563 ( .C1(n547), .C2(n546), .B(n545), .A(n544), .ZN(n3085) );
  nr02d0 U564 ( .A1(n549), .A2(n548), .ZN(n560) );
  nd02d0 U565 ( .A1(\hkspi/addr[5] ), .A2(n550), .ZN(n551) );
  nd02d0 U566 ( .A1(n556), .A2(n554), .ZN(n559) );
  nd02d0 U567 ( .A1(n555), .A2(\hkspi/addr[5] ), .ZN(n553) );
  oai211d1 U568 ( .C1(n560), .C2(n554), .A(n559), .B(n553), .ZN(n3084) );
  aon211d1 U569 ( .C1(n556), .C2(n558), .B(n555), .A(\hkspi/addr[6] ), .ZN(
        n557) );
  aon211d1 U570 ( .C1(n560), .C2(n559), .B(n558), .A(n557), .ZN(n3083) );
  aon211d1 U571 ( .C1(\hkspi/readmode ), .C2(n562), .B(rdstb), .A(n2316), .ZN(
        n561) );
  aoi21d1 U572 ( .B1(n563), .B2(n562), .A(n561), .ZN(n3082) );
  aoim21d1 U573 ( .B1(wrstb), .B2(\hkspi/writemode ), .A(n564), .ZN(n3081) );
  aoi22d1 U574 ( .A1(wbbd_busy), .A2(wbbd_data[0]), .B1(idata[0]), .B2(n2341), 
        .ZN(n1764) );
  inv0d1 U575 ( .I(n1764), .ZN(n3268) );
  nd02d0 U576 ( .A1(n817), .A2(n818), .ZN(n862) );
  inv0d0 U577 ( .I(n2264), .ZN(n2185) );
  nd02d0 U578 ( .A1(n2131), .A2(n1719), .ZN(n865) );
  nr02d0 U579 ( .A1(n2185), .A2(n865), .ZN(n565) );
  mx02d1 U580 ( .I0(hkspi_disable), .I1(n3268), .S(n565), .Z(n3080) );
  aoi211d1 U581 ( .C1(N867), .C2(N866), .A(N869), .B(N868), .ZN(n566) );
  nr04d0 U582 ( .A1(wb_adr_i[8]), .A2(wb_adr_i[9]), .A3(wb_adr_i[10]), .A4(
        wb_adr_i[11]), .ZN(n570) );
  nr04d0 U583 ( .A1(wb_adr_i[27]), .A2(wb_adr_i[12]), .A3(wb_adr_i[31]), .A4(
        wb_adr_i[28]), .ZN(n569) );
  nr04d0 U584 ( .A1(wb_adr_i[19]), .A2(wb_adr_i[14]), .A3(wb_adr_i[18]), .A4(
        wb_adr_i[17]), .ZN(n568) );
  inv0d0 U585 ( .I(wbbd_state[0]), .ZN(n808) );
  nd02d0 U586 ( .A1(n808), .A2(n581), .ZN(n3275) );
  inv0d0 U587 ( .I(n3275), .ZN(n3274) );
  oai211d1 U588 ( .C1(n579), .C2(n808), .A(wbbd_state[3]), .B(n3277), .ZN(n807) );
  oan211d1 U589 ( .C1(wrstb), .C2(rdstb), .B(n1718), .A(n797), .ZN(n574) );
  inv0d0 U590 ( .I(n574), .ZN(n578) );
  nd02d0 U591 ( .A1(n807), .A2(n578), .ZN(n582) );
  oan211d1 U592 ( .C1(n812), .C2(n803), .B(n3274), .A(n582), .ZN(n584) );
  nr03d1 U593 ( .A1(n3277), .A2(n579), .A3(n797), .ZN(n608) );
  inv0d0 U594 ( .I(n608), .ZN(n756) );
  nd02d0 U595 ( .A1(wbbd_state[3]), .A2(n807), .ZN(n802) );
  nd02d0 U596 ( .A1(n579), .A2(wbbd_state[3]), .ZN(n575) );
  oai211d1 U597 ( .C1(n584), .C2(n756), .A(n802), .B(n575), .ZN(n3079) );
  inv0d0 U598 ( .I(n582), .ZN(n577) );
  nr03d1 U599 ( .A1(n3277), .A2(n797), .A3(wbbd_state[1]), .ZN(n656) );
  inv0d0 U600 ( .I(n656), .ZN(n691) );
  inv0d0 U601 ( .I(n803), .ZN(n809) );
  nd02d0 U602 ( .A1(wbbd_state[0]), .A2(n809), .ZN(n576) );
  oai222d1 U603 ( .A1(n577), .A2(n691), .B1(n577), .B2(n576), .C1(n579), .C2(
        n582), .ZN(n3078) );
  nr03d1 U604 ( .A1(n579), .A2(n797), .A3(wbbd_state[2]), .ZN(n751) );
  inv0d0 U605 ( .I(n751), .ZN(n791) );
  oai21d1 U606 ( .B1(n579), .B2(n578), .A(wbbd_state[2]), .ZN(n580) );
  oai21d1 U607 ( .B1(n584), .B2(n791), .A(n580), .ZN(n3077) );
  oai21d1 U608 ( .B1(n809), .B2(n581), .A(n808), .ZN(n583) );
  oai22d1 U609 ( .A1(n584), .A2(n583), .B1(n808), .B2(n582), .ZN(n3076) );
  nr03d1 U610 ( .A1(n808), .A2(n803), .A3(wbbd_state[3]), .ZN(n726) );
  aoi22d1 U611 ( .A1(n726), .A2(wb_dat_i[0]), .B1(n751), .B2(wb_dat_i[8]), 
        .ZN(n589) );
  aoi22d1 U612 ( .A1(n656), .A2(wb_dat_i[16]), .B1(n608), .B2(wb_dat_i[24]), 
        .ZN(n588) );
  aoi22d1 U613 ( .A1(n656), .A2(wb_sel_i[2]), .B1(n608), .B2(wb_sel_i[3]), 
        .ZN(n586) );
  aoi22d1 U614 ( .A1(n726), .A2(wb_sel_i[0]), .B1(n751), .B2(wb_sel_i[1]), 
        .ZN(n585) );
  oaim21d1 U615 ( .B1(n586), .B2(n585), .A(wb_we_i), .ZN(n804) );
  nd02d0 U616 ( .A1(n804), .A2(wbbd_data[0]), .ZN(n587) );
  aon211d1 U617 ( .C1(n589), .C2(n588), .B(n804), .A(n587), .ZN(n3075) );
  aoi22d1 U618 ( .A1(n726), .A2(wb_dat_i[1]), .B1(n751), .B2(wb_dat_i[9]), 
        .ZN(n592) );
  aoi22d1 U619 ( .A1(n656), .A2(wb_dat_i[17]), .B1(n608), .B2(wb_dat_i[25]), 
        .ZN(n591) );
  nd02d0 U620 ( .A1(n804), .A2(wbbd_data[1]), .ZN(n590) );
  aon211d1 U621 ( .C1(n592), .C2(n591), .B(n804), .A(n590), .ZN(n3074) );
  aoi22d1 U622 ( .A1(n726), .A2(wb_dat_i[2]), .B1(n751), .B2(wb_dat_i[10]), 
        .ZN(n595) );
  aoi22d1 U623 ( .A1(n656), .A2(wb_dat_i[18]), .B1(n608), .B2(wb_dat_i[26]), 
        .ZN(n594) );
  nd02d0 U624 ( .A1(n804), .A2(wbbd_data[2]), .ZN(n593) );
  aon211d1 U625 ( .C1(n595), .C2(n594), .B(n804), .A(n593), .ZN(n3073) );
  aoi22d1 U626 ( .A1(n726), .A2(wb_dat_i[3]), .B1(n751), .B2(wb_dat_i[11]), 
        .ZN(n598) );
  aoi22d1 U627 ( .A1(n656), .A2(wb_dat_i[19]), .B1(n608), .B2(wb_dat_i[27]), 
        .ZN(n597) );
  nd02d0 U628 ( .A1(n804), .A2(wbbd_data[3]), .ZN(n596) );
  aon211d1 U629 ( .C1(n598), .C2(n597), .B(n804), .A(n596), .ZN(n3072) );
  aoi22d1 U630 ( .A1(n726), .A2(wb_dat_i[4]), .B1(n751), .B2(wb_dat_i[12]), 
        .ZN(n601) );
  aoi22d1 U631 ( .A1(n656), .A2(wb_dat_i[20]), .B1(n608), .B2(wb_dat_i[28]), 
        .ZN(n600) );
  nd02d0 U632 ( .A1(n804), .A2(wbbd_data[4]), .ZN(n599) );
  aon211d1 U633 ( .C1(n601), .C2(n600), .B(n804), .A(n599), .ZN(n3071) );
  aoi22d1 U634 ( .A1(n656), .A2(wb_dat_i[21]), .B1(n726), .B2(wb_dat_i[5]), 
        .ZN(n604) );
  aoi22d1 U635 ( .A1(n751), .A2(wb_dat_i[13]), .B1(n608), .B2(wb_dat_i[29]), 
        .ZN(n603) );
  nd02d0 U636 ( .A1(n804), .A2(wbbd_data[5]), .ZN(n602) );
  aon211d1 U637 ( .C1(n604), .C2(n603), .B(n804), .A(n602), .ZN(n3070) );
  aoi22d1 U638 ( .A1(n656), .A2(wb_dat_i[22]), .B1(n726), .B2(wb_dat_i[6]), 
        .ZN(n607) );
  aoi22d1 U639 ( .A1(n751), .A2(wb_dat_i[14]), .B1(n608), .B2(wb_dat_i[30]), 
        .ZN(n606) );
  nd02d0 U640 ( .A1(n804), .A2(wbbd_data[6]), .ZN(n605) );
  aon211d1 U641 ( .C1(n607), .C2(n606), .B(n804), .A(n605), .ZN(n3069) );
  aoi22d1 U642 ( .A1(n726), .A2(wb_dat_i[7]), .B1(n751), .B2(wb_dat_i[15]), 
        .ZN(n611) );
  aoi22d1 U643 ( .A1(n656), .A2(wb_dat_i[23]), .B1(n608), .B2(wb_dat_i[31]), 
        .ZN(n610) );
  nd02d0 U644 ( .A1(n804), .A2(wbbd_data[7]), .ZN(n609) );
  aon211d1 U645 ( .C1(n611), .C2(n610), .B(n804), .A(n609), .ZN(n3068) );
  inv0d1 U646 ( .I(N862), .ZN(n719) );
  inv0d0 U647 ( .I(N861), .ZN(n684) );
  nd02d0 U648 ( .A1(n719), .A2(n684), .ZN(n765) );
  inv0d0 U649 ( .I(n765), .ZN(n745) );
  inv0d0 U650 ( .I(N863), .ZN(n741) );
  nr03d0 U651 ( .A1(N867), .A2(N869), .A3(N868), .ZN(n627) );
  inv0d0 U652 ( .I(N866), .ZN(n631) );
  nd02d0 U653 ( .A1(n627), .A2(n631), .ZN(n612) );
  nr02d0 U654 ( .A1(N864), .A2(n612), .ZN(n766) );
  nd02d0 U655 ( .A1(n745), .A2(n712), .ZN(n742) );
  nr02d0 U656 ( .A1(N865), .A2(n612), .ZN(n615) );
  inv0d0 U657 ( .I(n778), .ZN(n669) );
  nd02d0 U658 ( .A1(N863), .A2(n669), .ZN(n787) );
  inv0d0 U659 ( .I(n787), .ZN(n784) );
  nr02d0 U660 ( .A1(n778), .A2(N863), .ZN(n673) );
  inv0d0 U661 ( .I(n673), .ZN(n767) );
  inv0d0 U662 ( .I(N860), .ZN(n665) );
  oai211d1 U663 ( .C1(n684), .C2(n665), .A(n673), .B(n719), .ZN(n613) );
  nr02d0 U664 ( .A1(n719), .A2(n731), .ZN(n717) );
  nd12d0 U665 ( .A1(n612), .A2(n632), .ZN(n629) );
  nd02d0 U666 ( .A1(n717), .A2(n722), .ZN(n650) );
  nd02d0 U667 ( .A1(n613), .A2(n650), .ZN(n718) );
  nr02d0 U668 ( .A1(n767), .A2(n718), .ZN(n624) );
  nr02d0 U669 ( .A1(N863), .A2(n699), .ZN(n782) );
  inv0d0 U670 ( .I(n786), .ZN(n639) );
  oai21d1 U671 ( .B1(n624), .B2(n782), .A(n639), .ZN(n614) );
  aon211d1 U672 ( .C1(n742), .C2(n736), .B(N860), .A(n614), .ZN(n753) );
  inv0d0 U673 ( .I(n782), .ZN(n744) );
  nr02d0 U674 ( .A1(N860), .A2(n684), .ZN(n685) );
  nd02d0 U675 ( .A1(N862), .A2(n685), .ZN(n759) );
  nd02d0 U676 ( .A1(n719), .A2(n685), .ZN(n618) );
  inv0d0 U677 ( .I(n618), .ZN(n701) );
  aon211d1 U678 ( .C1(N863), .C2(n615), .B(n712), .A(n701), .ZN(n616) );
  aon211d1 U679 ( .C1(n767), .C2(n744), .B(n759), .A(n616), .ZN(n667) );
  inv0d0 U680 ( .I(n759), .ZN(n670) );
  nd02d0 U681 ( .A1(n722), .A2(n670), .ZN(n617) );
  aon211d1 U682 ( .C1(n767), .C2(n744), .B(n618), .A(n617), .ZN(n679) );
  nd02d0 U683 ( .A1(n665), .A2(n745), .ZN(n700) );
  inv0d0 U684 ( .I(n700), .ZN(n635) );
  inv0d0 U685 ( .I(n722), .ZN(n758) );
  aoi21d1 U686 ( .B1(n758), .B2(n787), .A(n786), .ZN(n619) );
  oan211d1 U687 ( .C1(n673), .C2(n782), .B(n635), .A(n619), .ZN(n621) );
  oai211d1 U688 ( .C1(n787), .C2(n759), .A(n776), .B(n621), .ZN(n622) );
  nr04d0 U689 ( .A1(n753), .A2(n667), .A3(n679), .A4(n622), .ZN(n663) );
  nr02d0 U690 ( .A1(N861), .A2(n665), .ZN(n647) );
  nd02d0 U691 ( .A1(n647), .A2(n719), .ZN(n630) );
  nd02d0 U692 ( .A1(N862), .A2(n647), .ZN(n664) );
  or02d0 U693 ( .A1(n742), .A2(n665), .Z(n623) );
  nr02d0 U694 ( .A1(n630), .A2(n758), .ZN(n748) );
  inv0d0 U695 ( .I(n748), .ZN(n682) );
  oai211d1 U696 ( .C1(n664), .C2(n744), .A(n623), .B(n682), .ZN(n668) );
  nr02d0 U697 ( .A1(N862), .A2(n731), .ZN(n783) );
  nd02d0 U698 ( .A1(n783), .A2(n712), .ZN(n785) );
  inv0d0 U699 ( .I(n664), .ZN(n671) );
  nd02d0 U700 ( .A1(n712), .A2(n671), .ZN(n625) );
  inv0d0 U701 ( .I(n624), .ZN(n733) );
  nd02d0 U702 ( .A1(n671), .A2(n722), .ZN(n676) );
  aon211d1 U703 ( .C1(n758), .C2(n744), .B(n731), .A(n778), .ZN(n626) );
  nr04d0 U704 ( .A1(n680), .A2(n668), .A3(n763), .A4(n626), .ZN(n644) );
  inv0d0 U705 ( .I(n627), .ZN(n628) );
  nr04d0 U706 ( .A1(N864), .A2(N865), .A3(n628), .A4(n631), .ZN(n707) );
  nr02d0 U707 ( .A1(N863), .A2(n629), .ZN(n649) );
  nd02d0 U708 ( .A1(n649), .A2(n783), .ZN(n720) );
  nr02d0 U709 ( .A1(n647), .A2(n685), .ZN(n737) );
  nr02d0 U710 ( .A1(N862), .A2(n737), .ZN(n723) );
  inv0d0 U711 ( .I(n707), .ZN(n686) );
  nr02d0 U712 ( .A1(N863), .A2(n686), .ZN(n716) );
  oai21d1 U713 ( .B1(n723), .B2(n717), .A(n716), .ZN(n662) );
  aoi31d1 U714 ( .B1(n734), .B2(n720), .B3(n662), .A(n691), .ZN(n642) );
  inv0d0 U715 ( .I(n630), .ZN(n674) );
  nr04d0 U716 ( .A1(N863), .A2(N869), .A3(N868), .A4(n634), .ZN(n651) );
  nd02d0 U717 ( .A1(n649), .A2(n635), .ZN(n645) );
  inv0d0 U718 ( .I(n645), .ZN(n638) );
  inv0d0 U719 ( .I(n783), .ZN(n760) );
  nd02d0 U720 ( .A1(N863), .A2(n707), .ZN(n636) );
  oan211d1 U721 ( .C1(N861), .C2(N860), .B(n760), .A(n636), .ZN(n637) );
  aoi211d1 U722 ( .C1(n674), .C2(n651), .A(n638), .B(n637), .ZN(n743) );
  aoi21d1 U723 ( .B1(N861), .B2(N862), .A(n745), .ZN(n653) );
  nd02d0 U724 ( .A1(N860), .A2(n653), .ZN(n646) );
  an02d0 U725 ( .A1(n639), .A2(n651), .Z(n648) );
  aoi31d1 U726 ( .B1(n716), .B2(n700), .B3(n646), .A(n648), .ZN(n640) );
  oai21d1 U727 ( .B1(n783), .B2(n639), .A(n649), .ZN(n800) );
  inv0d0 U728 ( .I(n726), .ZN(n799) );
  aoi31d1 U729 ( .B1(n743), .B2(n640), .B3(n800), .A(n799), .ZN(n641) );
  aoi211d1 U730 ( .C1(wbbd_addr[0]), .C2(n797), .A(n642), .B(n641), .ZN(n643)
         );
  aon211d1 U731 ( .C1(n663), .C2(n644), .B(n791), .A(n643), .ZN(n3067) );
  oan211d1 U732 ( .C1(N863), .C2(N865), .B(n766), .A(n669), .ZN(n710) );
  oai211d1 U733 ( .C1(n710), .C2(n646), .A(n645), .B(n682), .ZN(n660) );
  nd02d0 U734 ( .A1(n716), .A2(n701), .ZN(n675) );
  nd02d0 U735 ( .A1(n707), .A2(n647), .ZN(n740) );
  nr02d0 U736 ( .A1(n741), .A2(n719), .ZN(n779) );
  aoi21d1 U737 ( .B1(n649), .B2(n674), .A(n648), .ZN(n683) );
  nd02d0 U738 ( .A1(n683), .A2(n650), .ZN(n770) );
  nd02d0 U739 ( .A1(n651), .A2(n719), .ZN(n738) );
  oaim22d1 U740 ( .A1(N861), .A2(n738), .B1(n670), .B2(n716), .ZN(n655) );
  nr02d0 U741 ( .A1(n669), .A2(n782), .ZN(n652) );
  oan211d1 U742 ( .C1(n653), .C2(n652), .B(n742), .A(n665), .ZN(n654) );
  nr03d0 U743 ( .A1(n770), .A2(n655), .A3(n654), .ZN(n709) );
  aon211d1 U744 ( .C1(n675), .C2(n740), .B(n779), .A(n709), .ZN(n659) );
  inv0d0 U745 ( .I(n797), .ZN(n693) );
  nr03d0 U746 ( .A1(n3277), .A2(n797), .A3(n720), .ZN(n796) );
  aoi31d1 U747 ( .B1(n716), .B2(n656), .B3(n717), .A(n796), .ZN(n730) );
  aoi211d1 U748 ( .C1(n734), .C2(n675), .A(n797), .B(n3277), .ZN(n695) );
  nd02d0 U749 ( .A1(N863), .A2(n695), .ZN(n757) );
  oai211d1 U750 ( .C1(n693), .C2(n657), .A(n730), .B(n757), .ZN(n658) );
  oan211d1 U751 ( .C1(n660), .C2(n659), .B(n726), .A(n658), .ZN(n661) );
  aon211d1 U752 ( .C1(n663), .C2(n662), .B(n791), .A(n661), .ZN(n3066) );
  oai22d1 U753 ( .A1(n665), .A2(n736), .B1(n664), .B2(n733), .ZN(n666) );
  nr03d0 U754 ( .A1(n668), .A2(n667), .A3(n666), .ZN(n735) );
  nd02d0 U755 ( .A1(n669), .A2(n779), .ZN(n711) );
  oai21d1 U756 ( .B1(n671), .B2(n670), .A(n712), .ZN(n672) );
  oai211d1 U757 ( .C1(n737), .C2(n711), .A(n672), .B(n720), .ZN(n790) );
  nd02d0 U758 ( .A1(n674), .A2(n673), .ZN(n677) );
  nd02d0 U759 ( .A1(n716), .A2(n717), .ZN(n690) );
  nr04d0 U760 ( .A1(n680), .A2(n679), .A3(n790), .A4(n678), .ZN(n698) );
  nr02d0 U761 ( .A1(n719), .A2(N861), .ZN(n681) );
  inv0d0 U762 ( .I(n681), .ZN(n703) );
  nr02d0 U763 ( .A1(n731), .A2(n738), .ZN(n705) );
  nd02d0 U764 ( .A1(n682), .A2(n690), .ZN(n704) );
  aon211d1 U765 ( .C1(n699), .C2(n711), .B(N861), .A(n683), .ZN(n780) );
  oai22d1 U766 ( .A1(n685), .A2(n779), .B1(n719), .B2(n684), .ZN(n687) );
  oai22d1 U767 ( .A1(N861), .A2(n778), .B1(n687), .B2(n686), .ZN(n688) );
  nr04d0 U768 ( .A1(n705), .A2(n704), .A3(n780), .A4(n688), .ZN(n689) );
  oai211d1 U769 ( .C1(n758), .C2(n703), .A(n689), .B(n720), .ZN(n696) );
  oai22d1 U770 ( .A1(n693), .A2(n692), .B1(n691), .B2(n690), .ZN(n694) );
  aoi211d1 U771 ( .C1(n726), .C2(n696), .A(n695), .B(n694), .ZN(n697) );
  aon211d1 U772 ( .C1(n735), .C2(n698), .B(n791), .A(n697), .ZN(n3065) );
  an02d0 U773 ( .A1(n699), .A2(n787), .Z(n777) );
  aon211d1 U774 ( .C1(n777), .C2(n767), .B(n700), .A(n800), .ZN(n728) );
  nd02d0 U775 ( .A1(N863), .A2(n701), .ZN(n702) );
  aon211d1 U776 ( .C1(n760), .C2(n703), .B(n779), .A(n702), .ZN(n706) );
  aoi211d1 U777 ( .C1(n707), .C2(n706), .A(n705), .B(n704), .ZN(n708) );
  oai211d1 U778 ( .C1(n710), .C2(n759), .A(n709), .B(n708), .ZN(n727) );
  oan211d1 U779 ( .C1(n719), .C2(n744), .B(n711), .A(n731), .ZN(n714) );
  inv0d0 U780 ( .I(n712), .ZN(n788) );
  aoi221d1 U781 ( .B1(n788), .B2(n744), .C1(N860), .C2(N861), .A(N862), .ZN(
        n713) );
  nr02d0 U782 ( .A1(n714), .A2(n713), .ZN(n793) );
  inv0d0 U783 ( .I(n734), .ZN(n715) );
  aoi21d1 U784 ( .B1(n716), .B2(n717), .A(n715), .ZN(n755) );
  inv0d0 U785 ( .I(n717), .ZN(n764) );
  aoi31d1 U786 ( .B1(n784), .B2(n719), .B3(n731), .A(n718), .ZN(n721) );
  oai211d1 U787 ( .C1(n764), .C2(n767), .A(n721), .B(n720), .ZN(n762) );
  aoi21d1 U788 ( .B1(n723), .B2(n722), .A(n762), .ZN(n724) );
  aoi31d1 U789 ( .B1(n793), .B2(n755), .B3(n724), .A(n791), .ZN(n725) );
  oan211d1 U790 ( .C1(n728), .C2(n727), .B(n726), .A(n725), .ZN(n729) );
  oaim211d1 U791 ( .C1(n797), .C2(wbbd_addr[3]), .A(n730), .B(n729), .ZN(n3064) );
  or02d0 U792 ( .A1(n731), .A2(n744), .Z(n732) );
  oai21d1 U793 ( .B1(n745), .B2(n767), .A(n736), .ZN(n769) );
  inv0d0 U794 ( .I(n737), .ZN(n739) );
  oai22d1 U795 ( .A1(n741), .A2(n740), .B1(n739), .B2(n738), .ZN(n747) );
  oai211d1 U796 ( .C1(n745), .C2(n744), .A(n743), .B(n742), .ZN(n746) );
  oaim22d1 U797 ( .A1(n749), .A2(n799), .B1(n797), .B2(wbbd_addr[4]), .ZN(n750) );
  oan211d1 U798 ( .C1(n753), .C2(n752), .B(n751), .A(n750), .ZN(n754) );
  aon211d1 U799 ( .C1(n757), .C2(n756), .B(n755), .A(n754), .ZN(n3063) );
  aoi31d1 U800 ( .B1(n760), .B2(n786), .B3(n759), .A(n758), .ZN(n761) );
  nr03d0 U801 ( .A1(n763), .A2(n762), .A3(n761), .ZN(n775) );
  nd02d0 U802 ( .A1(n800), .A2(n767), .ZN(n768) );
  nr03d0 U803 ( .A1(n770), .A2(n769), .A3(n768), .ZN(n771) );
  aoi21d1 U804 ( .B1(n772), .B2(n771), .A(n799), .ZN(n773) );
  aoi211d1 U805 ( .C1(wbbd_addr[5]), .C2(n797), .A(n796), .B(n773), .ZN(n774)
         );
  aon211d1 U806 ( .C1(n776), .C2(n775), .B(n791), .A(n774), .ZN(n3062) );
  aoi31d1 U807 ( .B1(N860), .B2(n779), .B3(n778), .A(n777), .ZN(n781) );
  aoi21d1 U808 ( .B1(N861), .B2(n781), .A(n780), .ZN(n801) );
  aoi21d1 U809 ( .B1(n784), .B2(n783), .A(n782), .ZN(n794) );
  aon211d1 U810 ( .C1(n788), .C2(n787), .B(n786), .A(n785), .ZN(n789) );
  nr02d0 U811 ( .A1(n790), .A2(n789), .ZN(n792) );
  aoi31d1 U812 ( .B1(n794), .B2(n793), .B3(n792), .A(n791), .ZN(n795) );
  aoi211d1 U813 ( .C1(wbbd_addr[6]), .C2(n797), .A(n796), .B(n795), .ZN(n798)
         );
  aon211d1 U814 ( .C1(n801), .C2(n800), .B(n799), .A(n798), .ZN(n3061) );
  nr02d0 U815 ( .A1(n3275), .A2(n803), .ZN(n811) );
  aoim21d1 U816 ( .B1(n802), .B2(wbbd_busy), .A(n811), .ZN(n3060) );
  aon211d1 U817 ( .C1(wbbd_state[3]), .C2(n803), .B(n808), .A(wbbd_write), 
        .ZN(n805) );
  aon211d1 U818 ( .C1(n806), .C2(wbbd_state[1]), .B(n805), .A(n804), .ZN(n3059) );
  nd02d0 U819 ( .A1(n807), .A2(wb_ack_o), .ZN(n810) );
  nd03d0 U820 ( .A1(wbbd_state[3]), .A2(n809), .A3(n808), .ZN(n3278) );
  aon211d1 U821 ( .C1(n812), .C2(n811), .B(n810), .A(n3278), .ZN(n3057) );
  inv0d0 U822 ( .I(n819), .ZN(n2290) );
  nd02d0 U823 ( .A1(n813), .A2(n815), .ZN(n2277) );
  inv0d0 U824 ( .I(n2277), .ZN(n2220) );
  nd02d0 U825 ( .A1(n2290), .A2(n2220), .ZN(n2171) );
  or02d0 U826 ( .A1(n2171), .A2(n1705), .Z(n839) );
  buffd1 U827 ( .I(n839), .Z(n3169) );
  nr02d0 U828 ( .A1(n1877), .A2(n3169), .ZN(n1710) );
  aoi22d1 U829 ( .A1(wbbd_busy), .A2(wbbd_data[1]), .B1(idata[1]), .B2(n2341), 
        .ZN(n1767) );
  inv0d1 U830 ( .I(n1767), .ZN(n3266) );
  inv0d0 U831 ( .I(n3266), .ZN(n1714) );
  aoim22d1 U832 ( .A1(n1710), .A2(n1714), .B1(irq_2_inputsrc), .B2(n1710), .Z(
        n3056) );
  inv0d0 U833 ( .I(serial_xfer), .ZN(n821) );
  nd02d0 U834 ( .A1(n815), .A2(n814), .ZN(n2288) );
  inv0d0 U835 ( .I(n2288), .ZN(n2137) );
  nr02d0 U836 ( .A1(n816), .A2(n830), .ZN(n860) );
  nd02d0 U837 ( .A1(n860), .A2(n834), .ZN(n851) );
  or02d0 U838 ( .A1(n851), .A2(n867), .Z(n2235) );
  inv0d0 U839 ( .I(n2235), .ZN(n2142) );
  nr04d0 U840 ( .A1(n819), .A2(n2288), .A3(n2235), .A4(n3268), .ZN(n820) );
  oan211d1 U841 ( .C1(n1705), .C2(n821), .B(n827), .A(n820), .ZN(n3055) );
  or02d0 U842 ( .A1(n871), .A2(n825), .Z(n1863) );
  nr02d0 U843 ( .A1(n1863), .A2(n2054), .ZN(n2139) );
  nd02d0 U844 ( .A1(n2139), .A2(n1719), .ZN(n822) );
  aoi22d1 U845 ( .A1(wbbd_busy), .A2(wbbd_data[5]), .B1(idata[5]), .B2(n2341), 
        .ZN(n1779) );
  inv0d0 U846 ( .I(n1779), .ZN(n3237) );
  inv0d1 U847 ( .I(n3237), .ZN(n1701) );
  aoi22d1 U848 ( .A1(wbbd_busy), .A2(wbbd_data[4]), .B1(idata[4]), .B2(n2341), 
        .ZN(n841) );
  inv0d0 U849 ( .I(n841), .ZN(n3245) );
  inv0d1 U850 ( .I(n3245), .ZN(n1702) );
  aoim22d1 U851 ( .A1(n824), .A2(n1702), .B1(mgmt_gpio_data[36]), .B2(n824), 
        .Z(n3053) );
  aoi22d1 U852 ( .A1(wbbd_busy), .A2(wbbd_data[3]), .B1(idata[3]), .B2(n2341), 
        .ZN(n837) );
  inv0d0 U853 ( .I(n837), .ZN(n3247) );
  inv0d1 U854 ( .I(n3247), .ZN(n846) );
  aoim22d1 U855 ( .A1(n824), .A2(n846), .B1(mgmt_gpio_data[35]), .B2(n824), 
        .Z(n3052) );
  inv0d1 U856 ( .I(n849), .ZN(n3260) );
  inv0d0 U857 ( .I(n3260), .ZN(n1713) );
  aoim22d1 U858 ( .A1(n824), .A2(n1713), .B1(mgmt_gpio_out[34]), .B2(n824), 
        .Z(n3051) );
  inv0d1 U859 ( .I(n1767), .ZN(n3242) );
  inv0d0 U860 ( .I(n3242), .ZN(n1759) );
  aoi22d1 U861 ( .A1(n824), .A2(n475), .B1(n823), .B2(n822), .ZN(n3050) );
  inv0d1 U862 ( .I(n1764), .ZN(n3272) );
  inv0d1 U863 ( .I(n3272), .ZN(n847) );
  aoim22d1 U864 ( .A1(n824), .A2(n847), .B1(mgmt_gpio_data_32), .B2(n824), .Z(
        n3049) );
  or02d0 U865 ( .A1(n867), .A2(n825), .Z(n1790) );
  buffd1 U866 ( .I(n874), .Z(n1711) );
  nr02d1 U867 ( .A1(n1790), .A2(n1711), .ZN(n826) );
  aoi22d1 U868 ( .A1(wbbd_busy), .A2(wbbd_data[7]), .B1(idata[7]), .B2(n2341), 
        .ZN(n855) );
  aoim22d1 U869 ( .A1(n826), .A2(n855), .B1(mgmt_gpio_out[31]), .B2(n826), .Z(
        n3048) );
  aoi22d1 U870 ( .A1(wbbd_busy), .A2(wbbd_data[6]), .B1(idata[6]), .B2(n2341), 
        .ZN(n876) );
  aoim22d1 U871 ( .A1(n826), .A2(n876), .B1(mgmt_gpio_out[30]), .B2(n826), .Z(
        n3047) );
  aoim22d1 U872 ( .A1(n826), .A2(n863), .B1(mgmt_gpio_out[29]), .B2(n826), .Z(
        n3046) );
  aoim22d1 U873 ( .A1(n826), .A2(n841), .B1(mgmt_gpio_out[28]), .B2(n826), .Z(
        n3045) );
  aoim22d1 U874 ( .A1(n826), .A2(n837), .B1(mgmt_gpio_out[27]), .B2(n826), .Z(
        n3044) );
  inv0d1 U875 ( .I(n849), .ZN(n3157) );
  inv0d0 U876 ( .I(n3157), .ZN(n836) );
  aoim22d1 U877 ( .A1(n826), .A2(n836), .B1(mgmt_gpio_out[26]), .B2(n826), .Z(
        n3043) );
  inv0d1 U878 ( .I(n1767), .ZN(n3270) );
  aoim22d1 U879 ( .A1(n826), .A2(n1767), .B1(mgmt_gpio_out[25]), .B2(n826), 
        .Z(n3042) );
  inv0d1 U880 ( .I(n1764), .ZN(n3233) );
  inv0d1 U881 ( .I(n3233), .ZN(n3181) );
  aoim22d1 U882 ( .A1(n826), .A2(n3181), .B1(mgmt_gpio_out[24]), .B2(n826), 
        .Z(n3041) );
  aoi22d1 U883 ( .A1(n828), .A2(n1759), .B1(n2181), .B2(n827), .ZN(n3040) );
  inv0d0 U884 ( .I(n876), .ZN(n3236) );
  inv0d1 U885 ( .I(n3236), .ZN(n878) );
  aoim22d1 U886 ( .A1(n828), .A2(n878), .B1(serial_bb_data_2), .B2(n828), .Z(
        n3039) );
  aoim22d1 U887 ( .A1(n828), .A2(n841), .B1(serial_bb_clock), .B2(n828), .Z(
        n3037) );
  aoim22d1 U888 ( .A1(n828), .A2(n837), .B1(serial_bb_load), .B2(n828), .Z(
        n3036) );
  aoim22d1 U889 ( .A1(n828), .A2(n836), .B1(serial_bb_resetn), .B2(n828), .Z(
        n3035) );
  an02d0 U890 ( .A1(n830), .A2(n829), .Z(n835) );
  nd02d0 U891 ( .A1(n861), .A2(n835), .ZN(n831) );
  or02d0 U892 ( .A1(n862), .A2(n831), .Z(n2076) );
  buffd1 U893 ( .I(n865), .Z(n872) );
  nr02d0 U894 ( .A1(n2076), .A2(n872), .ZN(n3248) );
  aoim22d1 U895 ( .A1(n3248), .A2(n836), .B1(\gpio_configure[37][10] ), .B2(
        n3248), .Z(n3034) );
  inv0d0 U896 ( .I(\gpio_configure[37][9] ), .ZN(n1508) );
  inv0d0 U897 ( .I(n3248), .ZN(n3246) );
  aoi22d1 U898 ( .A1(n3248), .A2(n475), .B1(n1508), .B2(n3246), .ZN(n3033) );
  inv0d0 U899 ( .I(\gpio_configure[37][8] ), .ZN(n1480) );
  aoi22d1 U900 ( .A1(n3248), .A2(n1764), .B1(n1480), .B2(n3246), .ZN(n3032) );
  nr02d1 U901 ( .A1(n1863), .A2(n1711), .ZN(n3186) );
  inv0d0 U902 ( .I(n855), .ZN(n3235) );
  inv0d0 U903 ( .I(\gpio_configure[37][7] ), .ZN(n1450) );
  inv0d0 U904 ( .I(n3186), .ZN(n3185) );
  aoi22d1 U905 ( .A1(n3186), .A2(n1786), .B1(n1450), .B2(n3185), .ZN(n3031) );
  inv0d0 U906 ( .I(\gpio_configure[37][6] ), .ZN(n1418) );
  aoi22d1 U907 ( .A1(n3186), .A2(n1782), .B1(n1418), .B2(n3185), .ZN(n3030) );
  aoim22d1 U908 ( .A1(n3186), .A2(n863), .B1(\gpio_configure[37][5] ), .B2(
        n3186), .Z(n3029) );
  inv0d0 U909 ( .I(n841), .ZN(n3230) );
  inv0d1 U910 ( .I(n3230), .ZN(n1775) );
  inv0d0 U911 ( .I(\gpio_configure[37][4] ), .ZN(n1360) );
  aoi22d1 U912 ( .A1(n3186), .A2(n1775), .B1(n1360), .B2(n3185), .ZN(n3028) );
  inv0d0 U913 ( .I(n837), .ZN(n3231) );
  inv0d1 U914 ( .I(n3231), .ZN(n1772) );
  aoi22d1 U915 ( .A1(n3186), .A2(n1772), .B1(mgmt_gpio_oeb[37]), .B2(n3185), 
        .ZN(n3027) );
  inv0d0 U916 ( .I(\gpio_configure[37][2] ), .ZN(n1306) );
  aoi22d1 U917 ( .A1(n3186), .A2(n849), .B1(n1306), .B2(n3185), .ZN(n3026) );
  inv0d0 U918 ( .I(\gpio_configure[36][10] ), .ZN(n1542) );
  inv0d0 U919 ( .I(n3105), .ZN(n3104) );
  aoi22d1 U920 ( .A1(n3105), .A2(n873), .B1(n1542), .B2(n3104), .ZN(n3025) );
  inv0d0 U921 ( .I(n3270), .ZN(n842) );
  aoim22d1 U922 ( .A1(n3105), .A2(n842), .B1(\gpio_configure[36][9] ), .B2(
        n3105), .Z(n3024) );
  aoim22d1 U923 ( .A1(n3105), .A2(n3181), .B1(\gpio_configure[36][8] ), .B2(
        n3105), .Z(n3023) );
  nr02d1 U924 ( .A1(n2076), .A2(n1711), .ZN(n3250) );
  inv0d1 U925 ( .I(n3235), .ZN(n852) );
  aoim22d1 U926 ( .A1(n3250), .A2(n852), .B1(\gpio_configure[36][7] ), .B2(
        n3250), .Z(n3022) );
  aoim22d1 U927 ( .A1(n3250), .A2(n878), .B1(\gpio_configure[36][6] ), .B2(
        n3250), .Z(n3021) );
  aoim22d1 U928 ( .A1(n3250), .A2(n863), .B1(\gpio_configure[36][5] ), .B2(
        n3250), .Z(n3020) );
  aoim22d1 U929 ( .A1(n3250), .A2(n841), .B1(\gpio_configure[36][4] ), .B2(
        n3250), .Z(n3019) );
  inv0d0 U930 ( .I(n3250), .ZN(n3249) );
  aoi22d1 U931 ( .A1(n3250), .A2(n1772), .B1(mgmt_gpio_oeb[36]), .B2(n3249), 
        .ZN(n3018) );
  aoim22d1 U932 ( .A1(n3250), .A2(n836), .B1(\gpio_configure[36][2] ), .B2(
        n3250), .Z(n3017) );
  nr02d1 U933 ( .A1(n831), .A2(n867), .ZN(n2041) );
  inv0d0 U934 ( .I(n2041), .ZN(n2072) );
  nr02d0 U935 ( .A1(n2072), .A2(n872), .ZN(n3141) );
  inv0d0 U936 ( .I(\gpio_configure[35][12] ), .ZN(n1631) );
  inv0d0 U937 ( .I(n3141), .ZN(n3140) );
  aoi22d1 U938 ( .A1(n3141), .A2(n1775), .B1(n1631), .B2(n3140), .ZN(n3016) );
  aoim22d1 U939 ( .A1(n3141), .A2(n837), .B1(\gpio_configure[35][11] ), .B2(
        n3141), .Z(n3015) );
  inv0d0 U940 ( .I(\gpio_configure[35][9] ), .ZN(n1509) );
  aoi22d1 U941 ( .A1(n3141), .A2(n1759), .B1(n1509), .B2(n3140), .ZN(n3014) );
  aoim22d1 U942 ( .A1(n3141), .A2(n3181), .B1(\gpio_configure[35][8] ), .B2(
        n3141), .Z(n3013) );
  nr02d1 U943 ( .A1(n2262), .A2(n874), .ZN(n3107) );
  inv0d0 U944 ( .I(\gpio_configure[35][7] ), .ZN(n1449) );
  inv0d0 U945 ( .I(n3107), .ZN(n3106) );
  aoi22d1 U946 ( .A1(n3107), .A2(n1786), .B1(n1449), .B2(n3106), .ZN(n3012) );
  aoim22d1 U947 ( .A1(n3107), .A2(n878), .B1(\gpio_configure[35][6] ), .B2(
        n3107), .Z(n3011) );
  inv0d0 U948 ( .I(\gpio_configure[35][5] ), .ZN(n1390) );
  aoi22d1 U949 ( .A1(n3107), .A2(n1779), .B1(n1390), .B2(n3106), .ZN(n3010) );
  aoim22d1 U950 ( .A1(n3107), .A2(n841), .B1(\gpio_configure[35][4] ), .B2(
        n3107), .Z(n3009) );
  aoim22d1 U951 ( .A1(n3107), .A2(n837), .B1(\gpio_configure[35][3] ), .B2(
        n3107), .Z(n3008) );
  inv0d0 U952 ( .I(\gpio_configure[35][2] ), .ZN(n1303) );
  aoi22d1 U953 ( .A1(n3107), .A2(n849), .B1(n1303), .B2(n3106), .ZN(n3007) );
  or02d0 U954 ( .A1(n831), .A2(n871), .Z(n1815) );
  inv0d0 U955 ( .I(\gpio_configure[34][12] ), .ZN(n1629) );
  inv0d0 U956 ( .I(n3192), .ZN(n3191) );
  aoi22d1 U957 ( .A1(n3192), .A2(n1775), .B1(n1629), .B2(n3191), .ZN(n3006) );
  inv0d0 U958 ( .I(\gpio_configure[34][11] ), .ZN(n1569) );
  aoi22d1 U959 ( .A1(n3192), .A2(n837), .B1(n1569), .B2(n3191), .ZN(n3005) );
  inv0d0 U960 ( .I(\gpio_configure[34][9] ), .ZN(n1512) );
  aoi22d1 U961 ( .A1(n3192), .A2(n1759), .B1(n1512), .B2(n3191), .ZN(n3004) );
  inv0d0 U962 ( .I(\gpio_configure[34][8] ), .ZN(n1477) );
  aoi22d1 U963 ( .A1(n3192), .A2(n3181), .B1(n1477), .B2(n3191), .ZN(n3003) );
  inv0d0 U964 ( .I(\gpio_configure[34][7] ), .ZN(n1448) );
  inv0d0 U965 ( .I(n3143), .ZN(n3142) );
  aoi22d1 U966 ( .A1(n3143), .A2(n1786), .B1(n1448), .B2(n3142), .ZN(n3002) );
  inv0d0 U967 ( .I(\gpio_configure[34][6] ), .ZN(n1421) );
  aoi22d1 U968 ( .A1(n3143), .A2(n1782), .B1(n1421), .B2(n3142), .ZN(n3001) );
  inv0d0 U969 ( .I(\gpio_configure[34][5] ), .ZN(n1389) );
  aoi22d1 U970 ( .A1(n3143), .A2(n1779), .B1(n1389), .B2(n3142), .ZN(n3000) );
  inv0d0 U971 ( .I(\gpio_configure[34][4] ), .ZN(n1363) );
  aoi22d1 U972 ( .A1(n3143), .A2(n1775), .B1(n1363), .B2(n3142), .ZN(n2999) );
  inv0d0 U973 ( .I(\gpio_configure[34][3] ), .ZN(n1332) );
  aoi22d1 U974 ( .A1(n3143), .A2(n837), .B1(n1332), .B2(n3142), .ZN(n2998) );
  inv0d0 U975 ( .I(\gpio_configure[34][2] ), .ZN(n1302) );
  aoi22d1 U976 ( .A1(n3143), .A2(n873), .B1(n1302), .B2(n3142), .ZN(n2997) );
  or02d0 U977 ( .A1(n832), .A2(n861), .Z(n833) );
  nr02d1 U978 ( .A1(n862), .A2(n833), .ZN(n2254) );
  nd02d0 U979 ( .A1(n2137), .A2(n1719), .ZN(n2333) );
  nd02d0 U980 ( .A1(n2254), .A2(n3228), .ZN(n3255) );
  inv0d0 U981 ( .I(n3255), .ZN(n3256) );
  aoim22d1 U982 ( .A1(n3256), .A2(n1775), .B1(\gpio_configure[33][12] ), .B2(
        n3256), .Z(n2996) );
  aoim22d1 U983 ( .A1(n3256), .A2(n1772), .B1(\gpio_configure[33][11] ), .B2(
        n3256), .Z(n2995) );
  aoim22d1 U984 ( .A1(n3256), .A2(n842), .B1(\gpio_configure[33][9] ), .B2(
        n3256), .Z(n2994) );
  inv0d0 U985 ( .I(\gpio_configure[33][8] ), .ZN(n1479) );
  aoi22d1 U986 ( .A1(n3256), .A2(n3181), .B1(n1479), .B2(n3255), .ZN(n2993) );
  nr02d1 U987 ( .A1(n1815), .A2(n874), .ZN(n3194) );
  inv0d0 U988 ( .I(\gpio_configure[33][7] ), .ZN(n1447) );
  inv0d0 U989 ( .I(n3194), .ZN(n3193) );
  aoi22d1 U990 ( .A1(n3194), .A2(n852), .B1(n1447), .B2(n3193), .ZN(n2992) );
  aoim22d1 U991 ( .A1(n3194), .A2(n878), .B1(\gpio_configure[33][6] ), .B2(
        n3194), .Z(n2991) );
  inv0d0 U992 ( .I(\gpio_configure[33][5] ), .ZN(n1391) );
  aoi22d1 U993 ( .A1(n3194), .A2(n1779), .B1(n1391), .B2(n3193), .ZN(n2990) );
  inv0d0 U994 ( .I(\gpio_configure[33][4] ), .ZN(n1359) );
  aoi22d1 U995 ( .A1(n3194), .A2(n841), .B1(n1359), .B2(n3193), .ZN(n2989) );
  inv0d0 U996 ( .I(\gpio_configure[33][3] ), .ZN(n1331) );
  aoi22d1 U997 ( .A1(n3194), .A2(n837), .B1(n1331), .B2(n3193), .ZN(n2988) );
  aoim22d1 U998 ( .A1(n3194), .A2(n836), .B1(\gpio_configure[33][2] ), .B2(
        n3194), .Z(n2987) );
  nr02d1 U999 ( .A1(n864), .A2(n833), .ZN(n2276) );
  nd02d0 U1000 ( .A1(n2276), .A2(n3228), .ZN(n3116) );
  inv0d0 U1001 ( .I(n3116), .ZN(n3117) );
  inv0d0 U1002 ( .I(\gpio_configure[32][12] ), .ZN(n1639) );
  aoi22d1 U1003 ( .A1(n3117), .A2(n841), .B1(n1639), .B2(n3116), .ZN(n2986) );
  inv0d0 U1004 ( .I(\gpio_configure[32][11] ), .ZN(n1568) );
  aoi22d1 U1005 ( .A1(n3117), .A2(n837), .B1(n1568), .B2(n3116), .ZN(n2985) );
  aoim22d1 U1006 ( .A1(n3117), .A2(n842), .B1(\gpio_configure[32][9] ), .B2(
        n3117), .Z(n2984) );
  inv0d0 U1007 ( .I(\gpio_configure[32][8] ), .ZN(n1481) );
  aoi22d1 U1008 ( .A1(n3117), .A2(n3181), .B1(n1481), .B2(n3116), .ZN(n2983)
         );
  aoim22d1 U1009 ( .A1(n3258), .A2(n852), .B1(\gpio_configure[32][7] ), .B2(
        n3258), .Z(n2982) );
  inv0d0 U1010 ( .I(\gpio_configure[32][6] ), .ZN(n1417) );
  aoi22d1 U1011 ( .A1(n3258), .A2(n1782), .B1(n1417), .B2(n3257), .ZN(n2981)
         );
  inv0d0 U1012 ( .I(\gpio_configure[32][5] ), .ZN(n1388) );
  aoi22d1 U1013 ( .A1(n3258), .A2(n1779), .B1(n1388), .B2(n3257), .ZN(n2980)
         );
  aoim22d1 U1014 ( .A1(n3258), .A2(n841), .B1(\gpio_configure[32][4] ), .B2(
        n3258), .Z(n2979) );
  inv0d0 U1015 ( .I(\gpio_configure[32][3] ), .ZN(n1333) );
  aoi22d1 U1016 ( .A1(n3258), .A2(n1772), .B1(n1333), .B2(n3257), .ZN(n2978)
         );
  aoim22d1 U1017 ( .A1(n3258), .A2(n836), .B1(\gpio_configure[32][2] ), .B2(
        n3258), .Z(n2977) );
  nr02d1 U1018 ( .A1(n833), .A2(n867), .ZN(n2258) );
  nd02d0 U1019 ( .A1(n2258), .A2(n3228), .ZN(n3152) );
  inv0d0 U1020 ( .I(n3152), .ZN(n3153) );
  aoim22d1 U1021 ( .A1(n3153), .A2(n841), .B1(\gpio_configure[31][12] ), .B2(
        n3153), .Z(n2976) );
  aoim22d1 U1022 ( .A1(n3153), .A2(n837), .B1(\gpio_configure[31][11] ), .B2(
        n3153), .Z(n2975) );
  aoim22d1 U1023 ( .A1(n3153), .A2(n842), .B1(\gpio_configure[31][9] ), .B2(
        n3153), .Z(n2974) );
  aoim22d1 U1024 ( .A1(n3153), .A2(n3181), .B1(\gpio_configure[31][8] ), .B2(
        n3153), .Z(n2973) );
  inv0d1 U1025 ( .I(n3118), .ZN(n3119) );
  aoim22d1 U1026 ( .A1(n3119), .A2(n852), .B1(\gpio_configure[31][7] ), .B2(
        n3119), .Z(n2972) );
  aoim22d1 U1027 ( .A1(n3119), .A2(n878), .B1(\gpio_configure[31][6] ), .B2(
        n3119), .Z(n2971) );
  aoim22d1 U1028 ( .A1(n3119), .A2(n863), .B1(\gpio_configure[31][5] ), .B2(
        n3119), .Z(n2970) );
  aoim22d1 U1029 ( .A1(n3119), .A2(n841), .B1(\gpio_configure[31][4] ), .B2(
        n3119), .Z(n2969) );
  aoim22d1 U1030 ( .A1(n3119), .A2(n837), .B1(\gpio_configure[31][3] ), .B2(
        n3119), .Z(n2968) );
  aoim22d1 U1031 ( .A1(n3119), .A2(n836), .B1(\gpio_configure[31][2] ), .B2(
        n3119), .Z(n2967) );
  nr02d1 U1032 ( .A1(n833), .A2(n871), .ZN(n2266) );
  nd02d0 U1033 ( .A1(n2266), .A2(n3228), .ZN(n3199) );
  inv0d0 U1034 ( .I(n3199), .ZN(n3200) );
  aoim22d1 U1035 ( .A1(n3200), .A2(n841), .B1(\gpio_configure[30][12] ), .B2(
        n3200), .Z(n2966) );
  aoim22d1 U1036 ( .A1(n3200), .A2(n1772), .B1(\gpio_configure[30][11] ), .B2(
        n3200), .Z(n2965) );
  aoim22d1 U1037 ( .A1(n3200), .A2(n842), .B1(\gpio_configure[30][9] ), .B2(
        n3200), .Z(n2964) );
  aoim22d1 U1038 ( .A1(n3200), .A2(n3181), .B1(\gpio_configure[30][8] ), .B2(
        n3200), .Z(n2963) );
  inv0d0 U1039 ( .I(n2258), .ZN(n1956) );
  nr02d1 U1040 ( .A1(n1956), .A2(n839), .ZN(n3155) );
  aoim22d1 U1041 ( .A1(n3155), .A2(n852), .B1(\gpio_configure[30][7] ), .B2(
        n3155), .Z(n2962) );
  aoim22d1 U1042 ( .A1(n3155), .A2(n878), .B1(\gpio_configure[30][6] ), .B2(
        n3155), .Z(n2961) );
  aoim22d1 U1043 ( .A1(n3155), .A2(n863), .B1(\gpio_configure[30][5] ), .B2(
        n3155), .Z(n2960) );
  aoim22d1 U1044 ( .A1(n3155), .A2(n1775), .B1(\gpio_configure[30][4] ), .B2(
        n3155), .Z(n2959) );
  aoim22d1 U1045 ( .A1(n3155), .A2(n837), .B1(\gpio_configure[30][3] ), .B2(
        n3155), .Z(n2958) );
  inv0d0 U1046 ( .I(\gpio_configure[30][2] ), .ZN(n1955) );
  inv0d0 U1047 ( .I(n3155), .ZN(n3154) );
  aoi22d1 U1048 ( .A1(n3155), .A2(n836), .B1(n1955), .B2(n3154), .ZN(n2957) );
  nd02d0 U1049 ( .A1(n835), .A2(n834), .ZN(n838) );
  nr02d1 U1050 ( .A1(n862), .A2(n838), .ZN(n2265) );
  nd02d0 U1051 ( .A1(n2265), .A2(n3228), .ZN(n3259) );
  inv0d0 U1052 ( .I(n3259), .ZN(n3261) );
  aoim22d1 U1053 ( .A1(n3261), .A2(n841), .B1(\gpio_configure[29][12] ), .B2(
        n3261), .Z(n2956) );
  aoim22d1 U1054 ( .A1(n3261), .A2(n837), .B1(\gpio_configure[29][11] ), .B2(
        n3261), .Z(n2955) );
  aoim22d1 U1055 ( .A1(n3261), .A2(n842), .B1(\gpio_configure[29][9] ), .B2(
        n3261), .Z(n2954) );
  aoim22d1 U1056 ( .A1(n3261), .A2(n3181), .B1(\gpio_configure[29][8] ), .B2(
        n3261), .Z(n2953) );
  nd12d0 U1057 ( .A1(n839), .A2(n2266), .ZN(n3201) );
  inv0d1 U1058 ( .I(n3201), .ZN(n3202) );
  aoim22d1 U1059 ( .A1(n3202), .A2(n852), .B1(\gpio_configure[29][7] ), .B2(
        n3202), .Z(n2952) );
  aoim22d1 U1060 ( .A1(n3202), .A2(n878), .B1(\gpio_configure[29][6] ), .B2(
        n3202), .Z(n2951) );
  aoim22d1 U1061 ( .A1(n3202), .A2(n863), .B1(\gpio_configure[29][5] ), .B2(
        n3202), .Z(n2950) );
  aoim22d1 U1062 ( .A1(n3202), .A2(n1775), .B1(\gpio_configure[29][4] ), .B2(
        n3202), .Z(n2949) );
  aoim22d1 U1063 ( .A1(n3202), .A2(n837), .B1(\gpio_configure[29][3] ), .B2(
        n3202), .Z(n2948) );
  aoim22d1 U1064 ( .A1(n3202), .A2(n836), .B1(\gpio_configure[29][2] ), .B2(
        n3202), .Z(n2947) );
  nr02d1 U1065 ( .A1(n864), .A2(n838), .ZN(n2253) );
  nd02d0 U1066 ( .A1(n2253), .A2(n3228), .ZN(n3120) );
  inv0d0 U1067 ( .I(n3120), .ZN(n3121) );
  aoim22d1 U1068 ( .A1(n3121), .A2(n841), .B1(\gpio_configure[28][12] ), .B2(
        n3121), .Z(n2946) );
  aoim22d1 U1069 ( .A1(n3121), .A2(n837), .B1(\gpio_configure[28][11] ), .B2(
        n3121), .Z(n2945) );
  aoim22d1 U1070 ( .A1(n3121), .A2(n842), .B1(\gpio_configure[28][9] ), .B2(
        n3121), .Z(n2944) );
  inv0d1 U1071 ( .I(n3272), .ZN(n868) );
  aoim22d1 U1072 ( .A1(n3121), .A2(n868), .B1(\gpio_configure[28][8] ), .B2(
        n3121), .Z(n2943) );
  nd12d0 U1073 ( .A1(n839), .A2(n2265), .ZN(n3262) );
  inv0d1 U1074 ( .I(n3262), .ZN(n3263) );
  aoim22d1 U1075 ( .A1(n3263), .A2(n852), .B1(\gpio_configure[28][7] ), .B2(
        n3263), .Z(n2942) );
  aoim22d1 U1076 ( .A1(n3263), .A2(n878), .B1(\gpio_configure[28][6] ), .B2(
        n3263), .Z(n2941) );
  aoim22d1 U1077 ( .A1(n3263), .A2(n863), .B1(\gpio_configure[28][5] ), .B2(
        n3263), .Z(n2940) );
  aoim22d1 U1078 ( .A1(n3263), .A2(n1775), .B1(\gpio_configure[28][4] ), .B2(
        n3263), .Z(n2939) );
  aoim22d1 U1079 ( .A1(n3263), .A2(n1772), .B1(\gpio_configure[28][3] ), .B2(
        n3263), .Z(n2938) );
  inv0d0 U1080 ( .I(n3157), .ZN(n840) );
  aoim22d1 U1081 ( .A1(n3263), .A2(n840), .B1(\gpio_configure[28][2] ), .B2(
        n3263), .Z(n2937) );
  nr02d1 U1082 ( .A1(n838), .A2(n867), .ZN(n2263) );
  nd02d0 U1083 ( .A1(n2263), .A2(n3228), .ZN(n3156) );
  inv0d0 U1084 ( .I(n3156), .ZN(n3158) );
  inv0d1 U1085 ( .I(n3245), .ZN(n866) );
  aoim22d1 U1086 ( .A1(n3158), .A2(n866), .B1(\gpio_configure[27][12] ), .B2(
        n3158), .Z(n2936) );
  aoim22d1 U1087 ( .A1(n3158), .A2(n1772), .B1(\gpio_configure[27][11] ), .B2(
        n3158), .Z(n2935) );
  aoim22d1 U1088 ( .A1(n3158), .A2(n842), .B1(\gpio_configure[27][9] ), .B2(
        n3158), .Z(n2934) );
  aoim22d1 U1089 ( .A1(n3158), .A2(n847), .B1(\gpio_configure[27][8] ), .B2(
        n3158), .Z(n2933) );
  nd12d0 U1090 ( .A1(n839), .A2(n2253), .ZN(n3122) );
  inv0d1 U1091 ( .I(n3122), .ZN(n3123) );
  aoim22d1 U1092 ( .A1(n3123), .A2(n852), .B1(\gpio_configure[27][7] ), .B2(
        n3123), .Z(n2932) );
  aoim22d1 U1093 ( .A1(n3123), .A2(n878), .B1(\gpio_configure[27][6] ), .B2(
        n3123), .Z(n2931) );
  aoim22d1 U1094 ( .A1(n3123), .A2(n863), .B1(\gpio_configure[27][5] ), .B2(
        n3123), .Z(n2930) );
  aoim22d1 U1095 ( .A1(n3123), .A2(n866), .B1(\gpio_configure[27][4] ), .B2(
        n3123), .Z(n2929) );
  inv0d1 U1096 ( .I(n3247), .ZN(n845) );
  aoim22d1 U1097 ( .A1(n3123), .A2(n845), .B1(\gpio_configure[27][3] ), .B2(
        n3123), .Z(n2928) );
  aoim22d1 U1098 ( .A1(n3123), .A2(n840), .B1(\gpio_configure[27][2] ), .B2(
        n3123), .Z(n2927) );
  nr02d1 U1099 ( .A1(n838), .A2(n871), .ZN(n2255) );
  nd02d0 U1100 ( .A1(n2255), .A2(n3228), .ZN(n3203) );
  inv0d0 U1101 ( .I(n3203), .ZN(n3205) );
  inv0d2 U1102 ( .I(n3245), .ZN(n856) );
  aoim22d1 U1103 ( .A1(n3205), .A2(n856), .B1(\gpio_configure[26][12] ), .B2(
        n3205), .Z(n2926) );
  aoim22d1 U1104 ( .A1(n3205), .A2(n845), .B1(\gpio_configure[26][11] ), .B2(
        n3205), .Z(n2925) );
  aoim22d1 U1105 ( .A1(n3205), .A2(n1767), .B1(\gpio_configure[26][9] ), .B2(
        n3205), .Z(n2924) );
  aoim22d1 U1106 ( .A1(n3205), .A2(n847), .B1(\gpio_configure[26][8] ), .B2(
        n3205), .Z(n2923) );
  nd12d0 U1107 ( .A1(n839), .A2(n2263), .ZN(n3159) );
  inv0d1 U1108 ( .I(n3159), .ZN(n3160) );
  aoim22d1 U1109 ( .A1(n3160), .A2(n852), .B1(\gpio_configure[26][7] ), .B2(
        n3160), .Z(n2922) );
  aoim22d1 U1110 ( .A1(n3160), .A2(n878), .B1(\gpio_configure[26][6] ), .B2(
        n3160), .Z(n2921) );
  aoim22d1 U1111 ( .A1(n3160), .A2(n863), .B1(\gpio_configure[26][5] ), .B2(
        n3160), .Z(n2920) );
  aoim22d1 U1112 ( .A1(n3160), .A2(n856), .B1(\gpio_configure[26][4] ), .B2(
        n3160), .Z(n2919) );
  aoim22d1 U1113 ( .A1(n3160), .A2(n845), .B1(\gpio_configure[26][3] ), .B2(
        n3160), .Z(n2918) );
  aoim22d1 U1114 ( .A1(n3160), .A2(n840), .B1(\gpio_configure[26][2] ), .B2(
        n3160), .Z(n2917) );
  nd02d0 U1115 ( .A1(n2264), .A2(n3228), .ZN(n3240) );
  inv0d0 U1116 ( .I(n3240), .ZN(n3241) );
  aoim22d1 U1117 ( .A1(n3241), .A2(n856), .B1(\gpio_configure[25][12] ), .B2(
        n3241), .Z(n2916) );
  aoim22d1 U1118 ( .A1(n3241), .A2(n845), .B1(\gpio_configure[25][11] ), .B2(
        n3241), .Z(n2915) );
  aoim22d1 U1119 ( .A1(n3241), .A2(n1767), .B1(\gpio_configure[25][9] ), .B2(
        n3241), .Z(n2914) );
  aoim22d1 U1120 ( .A1(n3241), .A2(n868), .B1(\gpio_configure[25][8] ), .B2(
        n3241), .Z(n2913) );
  inv0d1 U1121 ( .I(n3206), .ZN(n3207) );
  aoim22d1 U1122 ( .A1(n3207), .A2(n852), .B1(\gpio_configure[25][7] ), .B2(
        n3207), .Z(n2912) );
  aoim22d1 U1123 ( .A1(n3207), .A2(n878), .B1(\gpio_configure[25][6] ), .B2(
        n3207), .Z(n2911) );
  aoim22d1 U1124 ( .A1(n3207), .A2(n863), .B1(\gpio_configure[25][5] ), .B2(
        n3207), .Z(n2910) );
  aoim22d1 U1125 ( .A1(n3207), .A2(n1702), .B1(\gpio_configure[25][4] ), .B2(
        n3207), .Z(n2909) );
  aoim22d1 U1126 ( .A1(n3207), .A2(n845), .B1(\gpio_configure[25][3] ), .B2(
        n3207), .Z(n2908) );
  aoim22d1 U1127 ( .A1(n3207), .A2(n840), .B1(\gpio_configure[25][2] ), .B2(
        n3207), .Z(n2907) );
  nd02d0 U1128 ( .A1(n2195), .A2(n3228), .ZN(n3112) );
  inv0d0 U1129 ( .I(n3112), .ZN(n3113) );
  aoim22d1 U1130 ( .A1(n3113), .A2(n856), .B1(\gpio_configure[24][12] ), .B2(
        n3113), .Z(n2906) );
  aoim22d1 U1131 ( .A1(n3113), .A2(n845), .B1(\gpio_configure[24][11] ), .B2(
        n3113), .Z(n2905) );
  aoim22d1 U1132 ( .A1(n3113), .A2(n1767), .B1(\gpio_configure[24][9] ), .B2(
        n3113), .Z(n2904) );
  aoim22d1 U1133 ( .A1(n3113), .A2(n847), .B1(\gpio_configure[24][8] ), .B2(
        n3113), .Z(n2903) );
  nr02d1 U1134 ( .A1(n2185), .A2(n3169), .ZN(n3244) );
  aoim22d1 U1135 ( .A1(n3244), .A2(n855), .B1(\gpio_configure[24][7] ), .B2(
        n3244), .Z(n2902) );
  inv0d0 U1136 ( .I(\gpio_configure[24][6] ), .ZN(n2184) );
  inv0d0 U1137 ( .I(n3244), .ZN(n3243) );
  aoi22d1 U1138 ( .A1(n3244), .A2(n1782), .B1(n2184), .B2(n3243), .ZN(n2901)
         );
  aoim22d1 U1139 ( .A1(n3244), .A2(n863), .B1(\gpio_configure[24][5] ), .B2(
        n3244), .Z(n2900) );
  aoim22d1 U1140 ( .A1(n3244), .A2(n1702), .B1(\gpio_configure[24][4] ), .B2(
        n3244), .Z(n2899) );
  aoim22d1 U1141 ( .A1(n3244), .A2(n845), .B1(\gpio_configure[24][3] ), .B2(
        n3244), .Z(n2898) );
  aoim22d1 U1142 ( .A1(n3244), .A2(n840), .B1(\gpio_configure[24][2] ), .B2(
        n3244), .Z(n2897) );
  inv0d0 U1143 ( .I(n1790), .ZN(n2200) );
  nd02d0 U1144 ( .A1(n2200), .A2(n3228), .ZN(n3148) );
  inv0d0 U1145 ( .I(n3148), .ZN(n3149) );
  aoim22d1 U1146 ( .A1(n3149), .A2(n856), .B1(\gpio_configure[23][12] ), .B2(
        n3149), .Z(n2896) );
  aoim22d1 U1147 ( .A1(n3149), .A2(n845), .B1(\gpio_configure[23][11] ), .B2(
        n3149), .Z(n2895) );
  aoim22d1 U1148 ( .A1(n3149), .A2(n1767), .B1(\gpio_configure[23][9] ), .B2(
        n3149), .Z(n2894) );
  aoim22d1 U1149 ( .A1(n3149), .A2(n847), .B1(\gpio_configure[23][8] ), .B2(
        n3149), .Z(n2893) );
  nr02d1 U1150 ( .A1(n2093), .A2(n3169), .ZN(n3115) );
  aoim22d1 U1151 ( .A1(n3115), .A2(n852), .B1(\gpio_configure[23][7] ), .B2(
        n3115), .Z(n2892) );
  aoim22d1 U1152 ( .A1(n3115), .A2(n878), .B1(\gpio_configure[23][6] ), .B2(
        n3115), .Z(n2891) );
  aoim22d1 U1153 ( .A1(n3115), .A2(n863), .B1(\gpio_configure[23][5] ), .B2(
        n3115), .Z(n2890) );
  inv0d0 U1154 ( .I(\gpio_configure[23][4] ), .ZN(n2092) );
  inv0d0 U1155 ( .I(n3115), .ZN(n3114) );
  aoi22d1 U1156 ( .A1(n3115), .A2(n1775), .B1(n2092), .B2(n3114), .ZN(n2889)
         );
  aoim22d1 U1157 ( .A1(n3115), .A2(n845), .B1(\gpio_configure[23][3] ), .B2(
        n3115), .Z(n2888) );
  aoim22d1 U1158 ( .A1(n3115), .A2(n840), .B1(\gpio_configure[23][2] ), .B2(
        n3115), .Z(n2887) );
  inv0d0 U1159 ( .I(n1863), .ZN(n2001) );
  nd02d0 U1160 ( .A1(n2001), .A2(n3228), .ZN(n3187) );
  inv0d0 U1161 ( .I(n3187), .ZN(n3188) );
  aoim22d1 U1162 ( .A1(n3188), .A2(n856), .B1(\gpio_configure[22][12] ), .B2(
        n3188), .Z(n2886) );
  aoim22d1 U1163 ( .A1(n3188), .A2(n846), .B1(\gpio_configure[22][11] ), .B2(
        n3188), .Z(n2885) );
  aoim22d1 U1164 ( .A1(n3188), .A2(n1767), .B1(\gpio_configure[22][9] ), .B2(
        n3188), .Z(n2884) );
  aoim22d1 U1165 ( .A1(n3188), .A2(n868), .B1(\gpio_configure[22][8] ), .B2(
        n3188), .Z(n2883) );
  nr02d1 U1166 ( .A1(n1790), .A2(n3169), .ZN(n3151) );
  aoim22d1 U1167 ( .A1(n3151), .A2(n855), .B1(\gpio_configure[22][7] ), .B2(
        n3151), .Z(n2882) );
  aoim22d1 U1168 ( .A1(n3151), .A2(n878), .B1(\gpio_configure[22][6] ), .B2(
        n3151), .Z(n2881) );
  aoim22d1 U1169 ( .A1(n3151), .A2(n863), .B1(\gpio_configure[22][5] ), .B2(
        n3151), .Z(n2880) );
  aoim22d1 U1170 ( .A1(n3151), .A2(n856), .B1(\gpio_configure[22][4] ), .B2(
        n3151), .Z(n2879) );
  aoim22d1 U1171 ( .A1(n3151), .A2(n846), .B1(\gpio_configure[22][3] ), .B2(
        n3151), .Z(n2878) );
  aoim22d1 U1172 ( .A1(n3151), .A2(n840), .B1(\gpio_configure[22][2] ), .B2(
        n3151), .Z(n2877) );
  inv0d1 U1173 ( .I(n2076), .ZN(n2252) );
  nd02d0 U1174 ( .A1(n2252), .A2(n3228), .ZN(n3251) );
  inv0d0 U1175 ( .I(n3251), .ZN(n3252) );
  inv0d0 U1176 ( .I(\gpio_configure[21][12] ), .ZN(n2075) );
  aoi22d1 U1177 ( .A1(n3252), .A2(n841), .B1(n2075), .B2(n3251), .ZN(n2876) );
  aoim22d1 U1178 ( .A1(n3252), .A2(n846), .B1(\gpio_configure[21][11] ), .B2(
        n3252), .Z(n2875) );
  aoim22d1 U1179 ( .A1(n3252), .A2(n1767), .B1(\gpio_configure[21][9] ), .B2(
        n3252), .Z(n2874) );
  aoim22d1 U1180 ( .A1(n3252), .A2(n847), .B1(\gpio_configure[21][8] ), .B2(
        n3252), .Z(n2873) );
  nr02d1 U1181 ( .A1(n1863), .A2(n3169), .ZN(n3190) );
  aoim22d1 U1182 ( .A1(n3190), .A2(n855), .B1(\gpio_configure[21][7] ), .B2(
        n3190), .Z(n2872) );
  aoim22d1 U1183 ( .A1(n3190), .A2(n878), .B1(\gpio_configure[21][6] ), .B2(
        n3190), .Z(n2871) );
  aoim22d1 U1184 ( .A1(n3190), .A2(n863), .B1(\gpio_configure[21][5] ), .B2(
        n3190), .Z(n2870) );
  aoim22d1 U1185 ( .A1(n3190), .A2(n856), .B1(\gpio_configure[21][4] ), .B2(
        n3190), .Z(n2869) );
  aoim22d1 U1186 ( .A1(n3190), .A2(n846), .B1(\gpio_configure[21][3] ), .B2(
        n3190), .Z(n2868) );
  aoim22d1 U1187 ( .A1(n3190), .A2(n840), .B1(\gpio_configure[21][2] ), .B2(
        n3190), .Z(n2867) );
  inv0d1 U1188 ( .I(n2262), .ZN(n2225) );
  nd02d0 U1189 ( .A1(n2225), .A2(n3228), .ZN(n3108) );
  inv0d0 U1190 ( .I(n3108), .ZN(n3109) );
  aoim22d1 U1191 ( .A1(n3109), .A2(n856), .B1(\gpio_configure[20][12] ), .B2(
        n3109), .Z(n2866) );
  aoim22d1 U1192 ( .A1(n3109), .A2(n846), .B1(\gpio_configure[20][11] ), .B2(
        n3109), .Z(n2865) );
  aoim22d1 U1193 ( .A1(n3109), .A2(n1767), .B1(\gpio_configure[20][9] ), .B2(
        n3109), .Z(n2864) );
  aoim22d1 U1194 ( .A1(n3109), .A2(n868), .B1(\gpio_configure[20][8] ), .B2(
        n3109), .Z(n2863) );
  nr02d1 U1195 ( .A1(n2076), .A2(n3169), .ZN(n3254) );
  aoim22d1 U1196 ( .A1(n3254), .A2(n855), .B1(\gpio_configure[20][7] ), .B2(
        n3254), .Z(n2862) );
  aoim22d1 U1197 ( .A1(n3254), .A2(n876), .B1(\gpio_configure[20][6] ), .B2(
        n3254), .Z(n2861) );
  aoim22d1 U1198 ( .A1(n3254), .A2(n863), .B1(\gpio_configure[20][5] ), .B2(
        n3254), .Z(n2860) );
  aoim22d1 U1199 ( .A1(n3254), .A2(n856), .B1(\gpio_configure[20][4] ), .B2(
        n3254), .Z(n2859) );
  aoim22d1 U1200 ( .A1(n3254), .A2(n846), .B1(\gpio_configure[20][3] ), .B2(
        n3254), .Z(n2858) );
  aoim22d1 U1201 ( .A1(n3254), .A2(n840), .B1(\gpio_configure[20][2] ), .B2(
        n3254), .Z(n2857) );
  nd02d0 U1202 ( .A1(n2041), .A2(n3228), .ZN(n3144) );
  inv0d0 U1203 ( .I(n3144), .ZN(n3145) );
  inv0d0 U1204 ( .I(\gpio_configure[19][12] ), .ZN(n2071) );
  aoi22d1 U1205 ( .A1(n3145), .A2(n841), .B1(n2071), .B2(n3144), .ZN(n2856) );
  aoim22d1 U1206 ( .A1(n3145), .A2(n846), .B1(\gpio_configure[19][11] ), .B2(
        n3145), .Z(n2855) );
  inv0d0 U1207 ( .I(\gpio_configure[19][9] ), .ZN(n1875) );
  aoi22d1 U1208 ( .A1(n3145), .A2(n842), .B1(n1875), .B2(n3144), .ZN(n2854) );
  aoim22d1 U1209 ( .A1(n3145), .A2(n847), .B1(\gpio_configure[19][8] ), .B2(
        n3145), .Z(n2853) );
  nr02d1 U1210 ( .A1(n2262), .A2(n3169), .ZN(n3111) );
  inv0d0 U1211 ( .I(\gpio_configure[19][7] ), .ZN(n2261) );
  inv0d0 U1212 ( .I(n3111), .ZN(n3110) );
  aoi22d1 U1213 ( .A1(n3111), .A2(n852), .B1(n2261), .B2(n3110), .ZN(n2852) );
  aoim22d1 U1214 ( .A1(n3111), .A2(n876), .B1(\gpio_configure[19][6] ), .B2(
        n3111), .Z(n2851) );
  aoim22d1 U1215 ( .A1(n3111), .A2(n863), .B1(\gpio_configure[19][5] ), .B2(
        n3111), .Z(n2850) );
  aoim22d1 U1216 ( .A1(n3111), .A2(n856), .B1(\gpio_configure[19][4] ), .B2(
        n3111), .Z(n2849) );
  aoim22d1 U1217 ( .A1(n3111), .A2(n846), .B1(\gpio_configure[19][3] ), .B2(
        n3111), .Z(n2848) );
  inv0d1 U1218 ( .I(n849), .ZN(n3204) );
  inv0d1 U1219 ( .I(n3204), .ZN(n873) );
  aoim22d1 U1220 ( .A1(n3111), .A2(n873), .B1(\gpio_configure[19][2] ), .B2(
        n3111), .Z(n2847) );
  nd02d0 U1221 ( .A1(n2267), .A2(n3228), .ZN(n3195) );
  inv0d0 U1222 ( .I(n3195), .ZN(n3196) );
  aoim22d1 U1223 ( .A1(n3196), .A2(n856), .B1(\gpio_configure[18][12] ), .B2(
        n3196), .Z(n2846) );
  aoim22d1 U1224 ( .A1(n3196), .A2(n846), .B1(\gpio_configure[18][11] ), .B2(
        n3196), .Z(n2845) );
  inv0d0 U1225 ( .I(n3266), .ZN(n854) );
  aoim22d1 U1226 ( .A1(n3196), .A2(n854), .B1(\gpio_configure[18][9] ), .B2(
        n3196), .Z(n2844) );
  aoim22d1 U1227 ( .A1(n3196), .A2(n847), .B1(\gpio_configure[18][8] ), .B2(
        n3196), .Z(n2843) );
  nr02d1 U1228 ( .A1(n2072), .A2(n3169), .ZN(n3147) );
  aoim22d1 U1229 ( .A1(n3147), .A2(n1786), .B1(\gpio_configure[18][7] ), .B2(
        n3147), .Z(n2842) );
  aoim22d1 U1230 ( .A1(n3147), .A2(n878), .B1(\gpio_configure[18][6] ), .B2(
        n3147), .Z(n2841) );
  aoim22d1 U1231 ( .A1(n3147), .A2(n856), .B1(\gpio_configure[18][4] ), .B2(
        n3147), .Z(n2839) );
  aoim22d1 U1232 ( .A1(n3147), .A2(n845), .B1(\gpio_configure[18][3] ), .B2(
        n3147), .Z(n2838) );
  aoim22d1 U1233 ( .A1(n3147), .A2(n873), .B1(\gpio_configure[18][2] ), .B2(
        n3147), .Z(n2837) );
  or02d0 U1234 ( .A1(n843), .A2(n862), .Z(n2164) );
  nr02d1 U1235 ( .A1(n2164), .A2(n872), .ZN(n3217) );
  aoim22d1 U1236 ( .A1(n3217), .A2(n856), .B1(\gpio_configure[17][12] ), .B2(
        n3217), .Z(n2836) );
  aoim22d1 U1237 ( .A1(n3217), .A2(n846), .B1(\gpio_configure[17][11] ), .B2(
        n3217), .Z(n2835) );
  aoim22d1 U1238 ( .A1(n3217), .A2(n854), .B1(\gpio_configure[17][9] ), .B2(
        n3217), .Z(n2834) );
  aoim22d1 U1239 ( .A1(n3217), .A2(n847), .B1(\gpio_configure[17][8] ), .B2(
        n3217), .Z(n2833) );
  nr02d1 U1240 ( .A1(n1815), .A2(n3169), .ZN(n3198) );
  aoim22d1 U1241 ( .A1(n3198), .A2(n855), .B1(\gpio_configure[17][7] ), .B2(
        n3198), .Z(n2832) );
  aoim22d1 U1242 ( .A1(n3198), .A2(n876), .B1(\gpio_configure[17][6] ), .B2(
        n3198), .Z(n2831) );
  aoim22d1 U1243 ( .A1(n3198), .A2(n856), .B1(\gpio_configure[17][4] ), .B2(
        n3198), .Z(n2829) );
  aoim22d1 U1244 ( .A1(n3198), .A2(n845), .B1(\gpio_configure[17][3] ), .B2(
        n3198), .Z(n2828) );
  aoim22d1 U1245 ( .A1(n3198), .A2(n849), .B1(\gpio_configure[17][2] ), .B2(
        n3198), .Z(n2827) );
  nr02d1 U1246 ( .A1(n1877), .A2(n865), .ZN(n2324) );
  aoim22d1 U1247 ( .A1(n2324), .A2(n856), .B1(\gpio_configure[16][12] ), .B2(
        n2324), .Z(n2826) );
  aoim22d1 U1248 ( .A1(n2324), .A2(n846), .B1(\gpio_configure[16][11] ), .B2(
        n2324), .Z(n2825) );
  aoim22d1 U1249 ( .A1(n2324), .A2(n854), .B1(\gpio_configure[16][9] ), .B2(
        n2324), .Z(n2824) );
  aoim22d1 U1250 ( .A1(n2324), .A2(n847), .B1(\gpio_configure[16][8] ), .B2(
        n2324), .Z(n2823) );
  nr02d1 U1251 ( .A1(n2164), .A2(n1711), .ZN(n3219) );
  aoim22d1 U1252 ( .A1(n3219), .A2(n855), .B1(\gpio_configure[16][7] ), .B2(
        n3219), .Z(n2822) );
  aoim22d1 U1253 ( .A1(n3219), .A2(n1782), .B1(\gpio_configure[16][6] ), .B2(
        n3219), .Z(n2821) );
  aoim22d1 U1254 ( .A1(n3219), .A2(n856), .B1(\gpio_configure[16][4] ), .B2(
        n3219), .Z(n2819) );
  aoim22d1 U1255 ( .A1(n3219), .A2(n845), .B1(\gpio_configure[16][3] ), .B2(
        n3219), .Z(n2818) );
  aoim22d1 U1256 ( .A1(n3219), .A2(n849), .B1(\gpio_configure[16][2] ), .B2(
        n3219), .Z(n2817) );
  inv0d0 U1257 ( .I(n844), .ZN(n1914) );
  nr02d1 U1258 ( .A1(n1914), .A2(n872), .ZN(n3137) );
  aoim22d1 U1259 ( .A1(n3137), .A2(n856), .B1(\gpio_configure[15][12] ), .B2(
        n3137), .Z(n2816) );
  aoim22d1 U1260 ( .A1(n3137), .A2(n846), .B1(\gpio_configure[15][11] ), .B2(
        n3137), .Z(n2815) );
  aoim22d1 U1261 ( .A1(n3137), .A2(n854), .B1(\gpio_configure[15][9] ), .B2(
        n3137), .Z(n2814) );
  aoim22d1 U1262 ( .A1(n3137), .A2(n847), .B1(\gpio_configure[15][8] ), .B2(
        n3137), .Z(n2813) );
  aoim22d1 U1263 ( .A1(n2326), .A2(n855), .B1(\gpio_configure[15][7] ), .B2(
        n2326), .Z(n2812) );
  aoim22d1 U1264 ( .A1(n2326), .A2(n1782), .B1(\gpio_configure[15][6] ), .B2(
        n2326), .Z(n2811) );
  aoim22d1 U1265 ( .A1(n2326), .A2(n856), .B1(\gpio_configure[15][4] ), .B2(
        n2326), .Z(n2809) );
  aoim22d1 U1266 ( .A1(n2326), .A2(n845), .B1(\gpio_configure[15][3] ), .B2(
        n2326), .Z(n2808) );
  nr02d0 U1267 ( .A1(n1898), .A2(n872), .ZN(n3162) );
  aoim22d1 U1268 ( .A1(n3162), .A2(n856), .B1(\gpio_configure[14][12] ), .B2(
        n3162), .Z(n2806) );
  aoim22d1 U1269 ( .A1(n3162), .A2(n846), .B1(\gpio_configure[14][11] ), .B2(
        n3162), .Z(n2805) );
  inv0d0 U1270 ( .I(\gpio_configure[14][9] ), .ZN(n1897) );
  inv0d0 U1271 ( .I(n3162), .ZN(n3161) );
  aoi22d1 U1272 ( .A1(n3162), .A2(n475), .B1(n1897), .B2(n3161), .ZN(n2804) );
  aoim22d1 U1273 ( .A1(n3162), .A2(n847), .B1(\gpio_configure[14][8] ), .B2(
        n3162), .Z(n2803) );
  nr02d1 U1274 ( .A1(n1914), .A2(n1711), .ZN(n3139) );
  aoim22d1 U1275 ( .A1(n3139), .A2(n855), .B1(\gpio_configure[14][7] ), .B2(
        n3139), .Z(n2802) );
  aoim22d1 U1276 ( .A1(n3139), .A2(n876), .B1(\gpio_configure[14][6] ), .B2(
        n3139), .Z(n2801) );
  aoim22d1 U1277 ( .A1(n3139), .A2(n856), .B1(\gpio_configure[14][4] ), .B2(
        n3139), .Z(n2799) );
  inv0d1 U1278 ( .I(n3247), .ZN(n859) );
  aoim22d1 U1279 ( .A1(n3139), .A2(n859), .B1(\gpio_configure[14][3] ), .B2(
        n3139), .Z(n2798) );
  aoim22d1 U1280 ( .A1(n3139), .A2(n849), .B1(\gpio_configure[14][2] ), .B2(
        n3139), .Z(n2797) );
  nr02d1 U1281 ( .A1(n862), .A2(n851), .ZN(n2240) );
  inv0d0 U1282 ( .I(n2240), .ZN(n848) );
  nr02d1 U1283 ( .A1(n848), .A2(n872), .ZN(n3213) );
  aoim22d1 U1284 ( .A1(n3213), .A2(n856), .B1(\gpio_configure[13][12] ), .B2(
        n3213), .Z(n2796) );
  aoim22d1 U1285 ( .A1(n3213), .A2(n859), .B1(\gpio_configure[13][11] ), .B2(
        n3213), .Z(n2795) );
  aoim22d1 U1286 ( .A1(n3213), .A2(n854), .B1(\gpio_configure[13][9] ), .B2(
        n3213), .Z(n2794) );
  aoim22d1 U1287 ( .A1(n3213), .A2(n847), .B1(\gpio_configure[13][8] ), .B2(
        n3213), .Z(n2793) );
  aoim22d1 U1288 ( .A1(n3164), .A2(n1786), .B1(\gpio_configure[13][7] ), .B2(
        n3164), .Z(n2792) );
  aoim22d1 U1289 ( .A1(n3164), .A2(n876), .B1(\gpio_configure[13][6] ), .B2(
        n3164), .Z(n2791) );
  aoim22d1 U1290 ( .A1(n3164), .A2(n1702), .B1(\gpio_configure[13][4] ), .B2(
        n3164), .Z(n2789) );
  aoim22d1 U1291 ( .A1(n3164), .A2(n859), .B1(\gpio_configure[13][3] ), .B2(
        n3164), .Z(n2788) );
  nr02d1 U1292 ( .A1(n864), .A2(n851), .ZN(n2224) );
  inv0d0 U1293 ( .I(n2224), .ZN(n850) );
  nr02d1 U1294 ( .A1(n850), .A2(n865), .ZN(n2339) );
  aoim22d1 U1295 ( .A1(n2339), .A2(n866), .B1(\gpio_configure[12][12] ), .B2(
        n2339), .Z(n2786) );
  aoim22d1 U1296 ( .A1(n2339), .A2(n859), .B1(\gpio_configure[12][11] ), .B2(
        n2339), .Z(n2785) );
  aoim22d1 U1297 ( .A1(n2339), .A2(n854), .B1(\gpio_configure[12][9] ), .B2(
        n2339), .Z(n2784) );
  aoim22d1 U1298 ( .A1(n2339), .A2(n847), .B1(\gpio_configure[12][8] ), .B2(
        n2339), .Z(n2783) );
  nr02d1 U1299 ( .A1(n848), .A2(n1711), .ZN(n3215) );
  aoim22d1 U1300 ( .A1(n3215), .A2(n855), .B1(\gpio_configure[12][7] ), .B2(
        n3215), .Z(n2782) );
  aoim22d1 U1301 ( .A1(n3215), .A2(n1782), .B1(\gpio_configure[12][6] ), .B2(
        n3215), .Z(n2781) );
  aoim22d1 U1302 ( .A1(n3215), .A2(n1702), .B1(\gpio_configure[12][4] ), .B2(
        n3215), .Z(n2779) );
  aoim22d1 U1303 ( .A1(n3215), .A2(n859), .B1(\gpio_configure[12][3] ), .B2(
        n3215), .Z(n2778) );
  aoim22d1 U1304 ( .A1(n3215), .A2(n849), .B1(\gpio_configure[12][2] ), .B2(
        n3215), .Z(n2777) );
  nr02d1 U1305 ( .A1(n2235), .A2(n865), .ZN(n3125) );
  aoim22d1 U1306 ( .A1(n3125), .A2(n866), .B1(\gpio_configure[11][12] ), .B2(
        n3125), .Z(n2776) );
  aoim22d1 U1307 ( .A1(n3125), .A2(n859), .B1(\gpio_configure[11][11] ), .B2(
        n3125), .Z(n2775) );
  aoim22d1 U1308 ( .A1(n3125), .A2(n854), .B1(\gpio_configure[11][9] ), .B2(
        n3125), .Z(n2774) );
  aoim22d1 U1309 ( .A1(n3125), .A2(n868), .B1(\gpio_configure[11][8] ), .B2(
        n3125), .Z(n2773) );
  nr02d1 U1310 ( .A1(n850), .A2(n1711), .ZN(n2535) );
  aoim22d1 U1311 ( .A1(n2535), .A2(n855), .B1(\gpio_configure[11][7] ), .B2(
        n2535), .Z(n2772) );
  aoim22d1 U1312 ( .A1(n2535), .A2(n1782), .B1(\gpio_configure[11][6] ), .B2(
        n2535), .Z(n2771) );
  aoim22d1 U1313 ( .A1(n2535), .A2(n1702), .B1(\gpio_configure[11][4] ), .B2(
        n2535), .Z(n2769) );
  aoim22d1 U1314 ( .A1(n2535), .A2(n859), .B1(\gpio_configure[11][3] ), .B2(
        n2535), .Z(n2768) );
  aoim22d1 U1315 ( .A1(n2535), .A2(n873), .B1(\gpio_configure[11][2] ), .B2(
        n2535), .Z(n2767) );
  nr02d0 U1316 ( .A1(n871), .A2(n851), .ZN(n2067) );
  inv0d0 U1317 ( .I(n2067), .ZN(n3170) );
  nr02d1 U1318 ( .A1(n3170), .A2(n872), .ZN(n3166) );
  aoim22d1 U1319 ( .A1(n3166), .A2(n866), .B1(\gpio_configure[10][12] ), .B2(
        n3166), .Z(n2766) );
  aoim22d1 U1320 ( .A1(n3166), .A2(n859), .B1(\gpio_configure[10][11] ), .B2(
        n3166), .Z(n2765) );
  aoim22d1 U1321 ( .A1(n3166), .A2(n854), .B1(\gpio_configure[10][9] ), .B2(
        n3166), .Z(n2764) );
  aoim22d1 U1322 ( .A1(n3166), .A2(n868), .B1(\gpio_configure[10][8] ), .B2(
        n3166), .Z(n2763) );
  nr02d1 U1323 ( .A1(n2235), .A2(n874), .ZN(n3127) );
  inv0d0 U1324 ( .I(\gpio_configure[10][7] ), .ZN(n2234) );
  inv0d0 U1325 ( .I(n3127), .ZN(n3126) );
  aoi22d1 U1326 ( .A1(n3127), .A2(n852), .B1(n2234), .B2(n3126), .ZN(n2762) );
  aoim22d1 U1327 ( .A1(n3127), .A2(n1782), .B1(\gpio_configure[10][6] ), .B2(
        n3127), .Z(n2761) );
  aoim22d1 U1328 ( .A1(n3127), .A2(n1702), .B1(\gpio_configure[10][4] ), .B2(
        n3127), .Z(n2759) );
  aoim22d1 U1329 ( .A1(n3127), .A2(n859), .B1(\gpio_configure[10][3] ), .B2(
        n3127), .Z(n2758) );
  aoim22d1 U1330 ( .A1(n3127), .A2(n873), .B1(\gpio_configure[10][2] ), .B2(
        n3127), .Z(n2757) );
  nd02d0 U1331 ( .A1(n861), .A2(n853), .ZN(n857) );
  nr02d1 U1332 ( .A1(n862), .A2(n857), .ZN(n2282) );
  inv0d0 U1333 ( .I(n2282), .ZN(n1791) );
  nr02d1 U1334 ( .A1(n1791), .A2(n872), .ZN(n3225) );
  aoim22d1 U1335 ( .A1(n3225), .A2(n866), .B1(\gpio_configure[9][12] ), .B2(
        n3225), .Z(n2756) );
  aoim22d1 U1336 ( .A1(n3225), .A2(n859), .B1(\gpio_configure[9][11] ), .B2(
        n3225), .Z(n2755) );
  aoim22d1 U1337 ( .A1(n3225), .A2(n854), .B1(\gpio_configure[9][9] ), .B2(
        n3225), .Z(n2754) );
  aoim22d1 U1338 ( .A1(n3225), .A2(n868), .B1(\gpio_configure[9][8] ), .B2(
        n3225), .Z(n2753) );
  nr02d1 U1339 ( .A1(n3170), .A2(n1711), .ZN(n3168) );
  aoim22d1 U1340 ( .A1(n3168), .A2(n855), .B1(\gpio_configure[9][7] ), .B2(
        n3168), .Z(n2752) );
  aoim22d1 U1341 ( .A1(n3168), .A2(n876), .B1(\gpio_configure[9][6] ), .B2(
        n3168), .Z(n2751) );
  aoim22d1 U1342 ( .A1(n3168), .A2(n1702), .B1(\gpio_configure[9][4] ), .B2(
        n3168), .Z(n2749) );
  inv0d1 U1343 ( .I(n3247), .ZN(n1712) );
  aoim22d1 U1344 ( .A1(n3168), .A2(n1712), .B1(\gpio_configure[9][3] ), .B2(
        n3168), .Z(n2748) );
  aoim22d1 U1345 ( .A1(n3168), .A2(n873), .B1(\gpio_configure[9][2] ), .B2(
        n3168), .Z(n2747) );
  nr02d0 U1346 ( .A1(n857), .A2(n864), .ZN(n2205) );
  buffd1 U1347 ( .I(n2205), .Z(n2281) );
  inv0d0 U1348 ( .I(n2281), .ZN(n2334) );
  nr02d0 U1349 ( .A1(n2334), .A2(n872), .ZN(n2330) );
  aoim22d1 U1350 ( .A1(n2330), .A2(n866), .B1(\gpio_configure[8][12] ), .B2(
        n2330), .Z(n2746) );
  aoim22d1 U1351 ( .A1(n2330), .A2(n859), .B1(\gpio_configure[8][11] ), .B2(
        n2330), .Z(n2745) );
  inv0d0 U1352 ( .I(\gpio_configure[8][9] ), .ZN(n1901) );
  inv0d0 U1353 ( .I(n2330), .ZN(n2329) );
  aoi22d1 U1354 ( .A1(n2330), .A2(n1759), .B1(n1901), .B2(n2329), .ZN(n2744)
         );
  aoim22d1 U1355 ( .A1(n2330), .A2(n868), .B1(\gpio_configure[8][8] ), .B2(
        n2330), .Z(n2743) );
  nr02d1 U1356 ( .A1(n1791), .A2(n874), .ZN(n3227) );
  aoim22d1 U1357 ( .A1(n3227), .A2(n1786), .B1(\gpio_configure[8][7] ), .B2(
        n3227), .Z(n2742) );
  aoim22d1 U1358 ( .A1(n3227), .A2(n876), .B1(\gpio_configure[8][6] ), .B2(
        n3227), .Z(n2741) );
  aoim22d1 U1359 ( .A1(n3227), .A2(n1701), .B1(\gpio_configure[8][5] ), .B2(
        n3227), .Z(n2740) );
  aoim22d1 U1360 ( .A1(n3227), .A2(n866), .B1(\gpio_configure[8][4] ), .B2(
        n3227), .Z(n2739) );
  aoim22d1 U1361 ( .A1(n3227), .A2(n859), .B1(\gpio_configure[8][3] ), .B2(
        n3227), .Z(n2738) );
  aoim22d1 U1362 ( .A1(n3227), .A2(n873), .B1(\gpio_configure[8][2] ), .B2(
        n3227), .Z(n2737) );
  nr02d1 U1363 ( .A1(n857), .A2(n867), .ZN(n2241) );
  inv0d0 U1364 ( .I(n2241), .ZN(n1707) );
  nr02d1 U1365 ( .A1(n1707), .A2(n872), .ZN(n3133) );
  aoim22d1 U1366 ( .A1(n3133), .A2(n866), .B1(\gpio_configure[7][12] ), .B2(
        n3133), .Z(n2736) );
  aoim22d1 U1367 ( .A1(n3133), .A2(n1712), .B1(\gpio_configure[7][11] ), .B2(
        n3133), .Z(n2735) );
  aoim22d1 U1368 ( .A1(n3133), .A2(n1714), .B1(\gpio_configure[7][9] ), .B2(
        n3133), .Z(n2734) );
  aoim22d1 U1369 ( .A1(n3133), .A2(n868), .B1(\gpio_configure[7][8] ), .B2(
        n3133), .Z(n2733) );
  nr02d1 U1370 ( .A1(n2334), .A2(n1711), .ZN(n2332) );
  aoim22d1 U1371 ( .A1(n2332), .A2(n1786), .B1(\gpio_configure[7][7] ), .B2(
        n2332), .Z(n2732) );
  aoim22d1 U1372 ( .A1(n2332), .A2(n1782), .B1(\gpio_configure[7][6] ), .B2(
        n2332), .Z(n2731) );
  aoim22d1 U1373 ( .A1(n2332), .A2(n856), .B1(\gpio_configure[7][4] ), .B2(
        n2332), .Z(n2729) );
  aoim22d1 U1374 ( .A1(n2332), .A2(n859), .B1(\gpio_configure[7][3] ), .B2(
        n2332), .Z(n2728) );
  aoim22d1 U1375 ( .A1(n2332), .A2(n873), .B1(\gpio_configure[7][2] ), .B2(
        n2332), .Z(n2727) );
  nr02d1 U1376 ( .A1(n857), .A2(n871), .ZN(n858) );
  inv0d0 U1377 ( .I(n858), .ZN(n1703) );
  nr02d1 U1378 ( .A1(n1703), .A2(n872), .ZN(n3176) );
  aoim22d1 U1379 ( .A1(n3176), .A2(n866), .B1(\gpio_configure[6][12] ), .B2(
        n3176), .Z(n2726) );
  aoim22d1 U1380 ( .A1(n3176), .A2(n859), .B1(\gpio_configure[6][11] ), .B2(
        n3176), .Z(n2725) );
  aoim22d1 U1381 ( .A1(n3176), .A2(n1714), .B1(\gpio_configure[6][9] ), .B2(
        n3176), .Z(n2724) );
  aoim22d1 U1382 ( .A1(n3176), .A2(n868), .B1(\gpio_configure[6][8] ), .B2(
        n3176), .Z(n2723) );
  nr02d1 U1383 ( .A1(n1707), .A2(n874), .ZN(n3135) );
  aoim22d1 U1384 ( .A1(n3135), .A2(n1786), .B1(\gpio_configure[6][7] ), .B2(
        n3135), .Z(n2722) );
  aoim22d1 U1385 ( .A1(n3135), .A2(n1782), .B1(\gpio_configure[6][6] ), .B2(
        n3135), .Z(n2721) );
  aoim22d1 U1386 ( .A1(n3135), .A2(n866), .B1(\gpio_configure[6][4] ), .B2(
        n3135), .Z(n2719) );
  aoim22d1 U1387 ( .A1(n3135), .A2(n1712), .B1(\gpio_configure[6][3] ), .B2(
        n3135), .Z(n2718) );
  aoim22d1 U1388 ( .A1(n3135), .A2(n873), .B1(\gpio_configure[6][2] ), .B2(
        n3135), .Z(n2717) );
  nd02d0 U1389 ( .A1(n861), .A2(n860), .ZN(n870) );
  nr02d1 U1390 ( .A1(n862), .A2(n870), .ZN(n2222) );
  inv0d0 U1391 ( .I(n2222), .ZN(n1896) );
  aoim22d1 U1392 ( .A1(n3209), .A2(n866), .B1(\gpio_configure[5][12] ), .B2(
        n3209), .Z(n2716) );
  aoim22d1 U1393 ( .A1(n3209), .A2(n1712), .B1(\gpio_configure[5][11] ), .B2(
        n3209), .Z(n2715) );
  inv0d0 U1394 ( .I(\gpio_configure[5][9] ), .ZN(n1895) );
  inv0d0 U1395 ( .I(n3209), .ZN(n3208) );
  aoi22d1 U1396 ( .A1(n3209), .A2(n475), .B1(n1895), .B2(n3208), .ZN(n2714) );
  aoim22d1 U1397 ( .A1(n3209), .A2(n868), .B1(\gpio_configure[5][8] ), .B2(
        n3209), .Z(n2713) );
  nr02d1 U1398 ( .A1(n1703), .A2(n1711), .ZN(n3178) );
  aoim22d1 U1399 ( .A1(n3178), .A2(n1786), .B1(\gpio_configure[5][7] ), .B2(
        n3178), .Z(n2712) );
  aoim22d1 U1400 ( .A1(n3178), .A2(n876), .B1(\gpio_configure[5][6] ), .B2(
        n3178), .Z(n2711) );
  aoim22d1 U1401 ( .A1(n3178), .A2(n863), .B1(\gpio_configure[5][5] ), .B2(
        n3178), .Z(n2710) );
  aoim22d1 U1402 ( .A1(n3178), .A2(n866), .B1(\gpio_configure[5][4] ), .B2(
        n3178), .Z(n2709) );
  aoim22d1 U1403 ( .A1(n3178), .A2(n1712), .B1(\gpio_configure[5][3] ), .B2(
        n3178), .Z(n2708) );
  aoim22d1 U1404 ( .A1(n3178), .A2(n873), .B1(\gpio_configure[5][2] ), .B2(
        n3178), .Z(n2707) );
  nr02d1 U1405 ( .A1(n864), .A2(n870), .ZN(n2230) );
  inv0d0 U1406 ( .I(n2230), .ZN(n869) );
  nr02d1 U1407 ( .A1(n869), .A2(n865), .ZN(n2321) );
  aoim22d1 U1408 ( .A1(n2321), .A2(n866), .B1(\gpio_configure[4][12] ), .B2(
        n2321), .Z(n2706) );
  aoim22d1 U1409 ( .A1(n2321), .A2(n1712), .B1(\gpio_configure[4][11] ), .B2(
        n2321), .Z(n2705) );
  aoim22d1 U1410 ( .A1(n2321), .A2(n1714), .B1(\gpio_configure[4][9] ), .B2(
        n2321), .Z(n2704) );
  aoim22d1 U1411 ( .A1(n2321), .A2(n868), .B1(\gpio_configure[4][8] ), .B2(
        n2321), .Z(n2703) );
  nr02d1 U1412 ( .A1(n1896), .A2(n874), .ZN(n3211) );
  aoim22d1 U1413 ( .A1(n3211), .A2(n1786), .B1(\gpio_configure[4][7] ), .B2(
        n3211), .Z(n2702) );
  aoim22d1 U1414 ( .A1(n3211), .A2(n1782), .B1(\gpio_configure[4][6] ), .B2(
        n3211), .Z(n2701) );
  aoim22d1 U1415 ( .A1(n3211), .A2(n866), .B1(\gpio_configure[4][4] ), .B2(
        n3211), .Z(n2699) );
  aoim22d1 U1416 ( .A1(n3211), .A2(n1712), .B1(\gpio_configure[4][3] ), .B2(
        n3211), .Z(n2698) );
  aoim22d1 U1417 ( .A1(n3211), .A2(n873), .B1(\gpio_configure[4][2] ), .B2(
        n3211), .Z(n2697) );
  nr02d1 U1418 ( .A1(n867), .A2(n870), .ZN(n2238) );
  inv0d0 U1419 ( .I(n2238), .ZN(n2150) );
  nr02d1 U1420 ( .A1(n2150), .A2(n872), .ZN(n3131) );
  aoim22d1 U1421 ( .A1(n3131), .A2(n1702), .B1(\gpio_configure[3][12] ), .B2(
        n3131), .Z(n2696) );
  aoim22d1 U1422 ( .A1(n3131), .A2(n873), .B1(\gpio_configure[3][10] ), .B2(
        n3131), .Z(n2695) );
  aoim22d1 U1423 ( .A1(n3131), .A2(n1714), .B1(\gpio_configure[3][9] ), .B2(
        n3131), .Z(n2694) );
  aoim22d1 U1424 ( .A1(n3131), .A2(n868), .B1(\gpio_configure[3][8] ), .B2(
        n3131), .Z(n2693) );
  nr02d1 U1425 ( .A1(n869), .A2(n1711), .ZN(n3265) );
  aoim22d1 U1426 ( .A1(n3265), .A2(n1786), .B1(\gpio_configure[3][7] ), .B2(
        n3265), .Z(n2692) );
  aoim22d1 U1427 ( .A1(n3265), .A2(n1782), .B1(\gpio_configure[3][6] ), .B2(
        n3265), .Z(n2691) );
  aoim22d1 U1428 ( .A1(n3265), .A2(n1702), .B1(\gpio_configure[3][4] ), .B2(
        n3265), .Z(n2689) );
  aoim22d1 U1429 ( .A1(n3265), .A2(n1712), .B1(\gpio_configure[3][3] ), .B2(
        n3265), .Z(n2688) );
  aoim22d1 U1430 ( .A1(n3265), .A2(n1713), .B1(\gpio_configure[3][2] ), .B2(
        n3265), .Z(n2687) );
  aoim22d1 U1431 ( .A1(n3265), .A2(n1767), .B1(\gpio_configure[3][1] ), .B2(
        n3265), .Z(n2686) );
  nr02d1 U1432 ( .A1(n871), .A2(n870), .ZN(n2242) );
  inv0d0 U1433 ( .I(n2242), .ZN(n875) );
  nr02d1 U1434 ( .A1(n875), .A2(n872), .ZN(n3184) );
  aoim22d1 U1435 ( .A1(n3184), .A2(n1702), .B1(\gpio_configure[2][12] ), .B2(
        n3184), .Z(n2685) );
  aoim22d1 U1436 ( .A1(n3184), .A2(n1712), .B1(\gpio_configure[2][11] ), .B2(
        n3184), .Z(n2684) );
  aoim22d1 U1437 ( .A1(n3184), .A2(n1714), .B1(\gpio_configure[2][9] ), .B2(
        n3184), .Z(n2683) );
  aoim22d1 U1438 ( .A1(n3184), .A2(n1764), .B1(\gpio_configure[2][8] ), .B2(
        n3184), .Z(n2682) );
  nr02d1 U1439 ( .A1(n2150), .A2(n1711), .ZN(n3269) );
  aoim22d1 U1440 ( .A1(n3269), .A2(n1786), .B1(\gpio_configure[2][7] ), .B2(
        n3269), .Z(n2681) );
  aoim22d1 U1441 ( .A1(n3269), .A2(n876), .B1(\gpio_configure[2][6] ), .B2(
        n3269), .Z(n2680) );
  inv0d0 U1442 ( .I(\gpio_configure[2][5] ), .ZN(n2149) );
  inv0d0 U1443 ( .I(n3269), .ZN(n3267) );
  aoi22d1 U1444 ( .A1(n3269), .A2(n1779), .B1(n2149), .B2(n3267), .ZN(n2679)
         );
  aoim22d1 U1445 ( .A1(n3269), .A2(n1702), .B1(\gpio_configure[2][4] ), .B2(
        n3269), .Z(n2678) );
  aoim22d1 U1446 ( .A1(n3269), .A2(n1712), .B1(\gpio_configure[2][3] ), .B2(
        n3269), .Z(n2677) );
  aoim22d1 U1447 ( .A1(n3269), .A2(n1713), .B1(\gpio_configure[2][2] ), .B2(
        n3269), .Z(n2676) );
  inv0d2 U1448 ( .I(n2164), .ZN(n2256) );
  nd02d0 U1449 ( .A1(n2256), .A2(n3228), .ZN(n3220) );
  inv0d0 U1450 ( .I(n3220), .ZN(n3221) );
  aoim22d1 U1451 ( .A1(n3221), .A2(n873), .B1(\gpio_configure[1][10] ), .B2(
        n3221), .Z(n2675) );
  inv0d0 U1452 ( .I(\gpio_configure[1][9] ), .ZN(n1880) );
  aoi22d1 U1453 ( .A1(n3221), .A2(n475), .B1(n1880), .B2(n3220), .ZN(n2674) );
  aoim22d1 U1454 ( .A1(n3221), .A2(n1764), .B1(\gpio_configure[1][8] ), .B2(
        n3221), .Z(n2673) );
  nr02d1 U1455 ( .A1(n875), .A2(n874), .ZN(n3273) );
  aoim22d1 U1456 ( .A1(n3273), .A2(n1786), .B1(\gpio_configure[1][7] ), .B2(
        n3273), .Z(n2672) );
  aoim22d1 U1457 ( .A1(n3273), .A2(n876), .B1(\gpio_configure[1][6] ), .B2(
        n3273), .Z(n2671) );
  aoim22d1 U1458 ( .A1(n3273), .A2(n1702), .B1(\gpio_configure[1][4] ), .B2(
        n3273), .Z(n2669) );
  inv0d0 U1459 ( .I(n3273), .ZN(n3271) );
  aoi22d1 U1460 ( .A1(n3273), .A2(n1772), .B1(n877), .B2(n3271), .ZN(n2668) );
  aoim22d1 U1461 ( .A1(n3273), .A2(n1713), .B1(\gpio_configure[1][2] ), .B2(
        n3273), .Z(n2667) );
  nd02d0 U1462 ( .A1(n2223), .A2(n3228), .ZN(n2327) );
  inv0d0 U1463 ( .I(n2327), .ZN(n2328) );
  aoim22d1 U1464 ( .A1(n2328), .A2(n1713), .B1(\gpio_configure[0][10] ), .B2(
        n2328), .Z(n2666) );
  inv0d0 U1465 ( .I(\gpio_configure[0][9] ), .ZN(n1876) );
  aoi22d1 U1466 ( .A1(n2328), .A2(n1759), .B1(n1876), .B2(n2327), .ZN(n2665)
         );
  aoim22d1 U1467 ( .A1(n2328), .A2(n3181), .B1(\gpio_configure[0][8] ), .B2(
        n2328), .Z(n2664) );
  nr02d1 U1468 ( .A1(n2164), .A2(n3169), .ZN(n3223) );
  aoim22d1 U1469 ( .A1(n3223), .A2(n1786), .B1(\gpio_configure[0][7] ), .B2(
        n3223), .Z(n2663) );
  aoim22d1 U1470 ( .A1(n3223), .A2(n878), .B1(\gpio_configure[0][6] ), .B2(
        n3223), .Z(n2662) );
  inv0d0 U1471 ( .I(\gpio_configure[0][5] ), .ZN(n2163) );
  inv0d0 U1472 ( .I(n3223), .ZN(n3222) );
  aoi22d1 U1473 ( .A1(n3223), .A2(n1779), .B1(n2163), .B2(n3222), .ZN(n2661)
         );
  aoim22d1 U1474 ( .A1(n3223), .A2(n1702), .B1(\gpio_configure[0][4] ), .B2(
        n3223), .Z(n2660) );
  aoi22d1 U1475 ( .A1(n3223), .A2(n1772), .B1(n879), .B2(n3222), .ZN(n2659) );
  aoim22d1 U1476 ( .A1(n3223), .A2(n1713), .B1(\gpio_configure[0][2] ), .B2(
        n3223), .Z(n2658) );
  inv0d0 U1477 ( .I(pad_count_1[1]), .ZN(n881) );
  inv0d0 U1478 ( .I(pad_count_1[0]), .ZN(n1686) );
  nd02d0 U1479 ( .A1(n881), .A2(n1686), .ZN(n1688) );
  nr02d0 U1480 ( .A1(n1688), .A2(pad_count_1[2]), .ZN(n1690) );
  inv0d0 U1481 ( .I(n1690), .ZN(n1693) );
  nd02d0 U1482 ( .A1(pad_count_1[4]), .A2(pad_count_1[3]), .ZN(n880) );
  nr02d1 U1483 ( .A1(n1693), .A2(n880), .ZN(n1161) );
  nd02d0 U1484 ( .A1(pad_count_1[0]), .A2(n881), .ZN(n905) );
  inv0d0 U1485 ( .I(pad_count_1[3]), .ZN(n1694) );
  nr02d0 U1486 ( .A1(pad_count_1[4]), .A2(n1694), .ZN(n1698) );
  inv0d0 U1487 ( .I(pad_count_1[2]), .ZN(n1691) );
  nd02d0 U1488 ( .A1(n1698), .A2(n1691), .ZN(n900) );
  nr02d1 U1489 ( .A1(n905), .A2(n900), .ZN(n1186) );
  aoi22d1 U1490 ( .A1(\gpio_configure[24][12] ), .A2(n1161), .B1(
        \gpio_configure[9][12] ), .B2(n1186), .ZN(n886) );
  nd02d0 U1491 ( .A1(pad_count_1[1]), .A2(pad_count_1[0]), .ZN(n903) );
  nr02d0 U1492 ( .A1(pad_count_1[4]), .A2(pad_count_1[3]), .ZN(n882) );
  nd02d0 U1493 ( .A1(n882), .A2(n1691), .ZN(n892) );
  nr02d1 U1494 ( .A1(n903), .A2(n892), .ZN(n1162) );
  nd02d0 U1495 ( .A1(pad_count_1[2]), .A2(n882), .ZN(n904) );
  nr02d1 U1496 ( .A1(n903), .A2(n904), .ZN(n1173) );
  aoi22d1 U1497 ( .A1(\gpio_configure[3][12] ), .A2(n1162), .B1(
        \gpio_configure[7][12] ), .B2(n1173), .ZN(n885) );
  nd03d0 U1498 ( .A1(pad_count_1[2]), .A2(pad_count_1[4]), .A3(pad_count_1[3]), 
        .ZN(n902) );
  nr02d1 U1499 ( .A1(n905), .A2(n902), .ZN(n1203) );
  nr02d1 U1500 ( .A1(n905), .A2(n892), .ZN(n1202) );
  aoi22d1 U1501 ( .A1(\gpio_configure[29][12] ), .A2(n1203), .B1(
        \gpio_configure[1][12] ), .B2(n1202), .ZN(n884) );
  nd02d0 U1502 ( .A1(pad_count_1[1]), .A2(n1686), .ZN(n899) );
  nd03d0 U1503 ( .A1(pad_count_1[4]), .A2(n1691), .A3(n1694), .ZN(n901) );
  nr02d1 U1504 ( .A1(n899), .A2(n901), .ZN(n1177) );
  an03d1 U1505 ( .A1(n1694), .A2(pad_count_1[4]), .A3(n1690), .Z(n1697) );
  aoi22d1 U1506 ( .A1(\gpio_configure[18][12] ), .A2(n1177), .B1(
        \gpio_configure[16][12] ), .B2(n1697), .ZN(n883) );
  nd03d0 U1507 ( .A1(pad_count_1[4]), .A2(pad_count_1[2]), .A3(n1694), .ZN(
        n897) );
  nr02d1 U1508 ( .A1(n899), .A2(n897), .ZN(n1200) );
  nr02d1 U1509 ( .A1(n904), .A2(n899), .ZN(n1176) );
  aoi22d1 U1510 ( .A1(\gpio_configure[22][12] ), .A2(n1200), .B1(
        \gpio_configure[6][12] ), .B2(n1176), .ZN(n890) );
  an02d1 U1511 ( .A1(n1698), .A2(n1690), .Z(n1167) );
  nr02d1 U1512 ( .A1(n1688), .A2(n904), .ZN(n1189) );
  aoi22d1 U1513 ( .A1(\gpio_configure[8][12] ), .A2(n1167), .B1(
        \gpio_configure[4][12] ), .B2(n1189), .ZN(n889) );
  nd02d0 U1514 ( .A1(pad_count_1[2]), .A2(n1698), .ZN(n891) );
  nr02d1 U1515 ( .A1(n905), .A2(n891), .ZN(n1187) );
  nr02d1 U1516 ( .A1(n903), .A2(n891), .ZN(n1188) );
  aoi22d1 U1517 ( .A1(\gpio_configure[13][12] ), .A2(n1187), .B1(
        \gpio_configure[15][12] ), .B2(n1188), .ZN(n888) );
  nr02d1 U1518 ( .A1(n1688), .A2(n897), .ZN(n1163) );
  nr02d1 U1519 ( .A1(n900), .A2(n903), .ZN(n1168) );
  aoi22d1 U1520 ( .A1(\gpio_configure[20][12] ), .A2(n1163), .B1(
        \gpio_configure[11][12] ), .B2(n1168), .ZN(n887) );
  nd03d0 U1521 ( .A1(pad_count_1[4]), .A2(pad_count_1[3]), .A3(n1691), .ZN(
        n898) );
  nr02d1 U1522 ( .A1(n899), .A2(n898), .ZN(n1179) );
  nr02d1 U1523 ( .A1(n902), .A2(n899), .ZN(n1164) );
  aoi22d1 U1524 ( .A1(\gpio_configure[26][12] ), .A2(n1179), .B1(
        \gpio_configure[30][12] ), .B2(n1164), .ZN(n896) );
  nr02d1 U1525 ( .A1(n905), .A2(n898), .ZN(n1201) );
  nr02d1 U1526 ( .A1(n1688), .A2(n902), .ZN(n1165) );
  aoi22d1 U1527 ( .A1(\gpio_configure[25][12] ), .A2(n1201), .B1(
        \gpio_configure[28][12] ), .B2(n1165), .ZN(n895) );
  nr02d1 U1528 ( .A1(n899), .A2(n891), .ZN(n1197) );
  nr02d1 U1529 ( .A1(n1688), .A2(n891), .ZN(n1180) );
  aoi22d1 U1530 ( .A1(\gpio_configure[14][12] ), .A2(n1197), .B1(
        \gpio_configure[12][12] ), .B2(n1180), .ZN(n894) );
  nr02d1 U1531 ( .A1(n903), .A2(n897), .ZN(n1190) );
  nr02d1 U1532 ( .A1(n892), .A2(n899), .ZN(n1178) );
  aoi22d1 U1533 ( .A1(\gpio_configure[23][12] ), .A2(n1190), .B1(
        \gpio_configure[2][12] ), .B2(n1178), .ZN(n893) );
  nr02d1 U1534 ( .A1(n905), .A2(n897), .ZN(n1196) );
  nr02d1 U1535 ( .A1(n903), .A2(n898), .ZN(n1198) );
  aoi22d1 U1536 ( .A1(\gpio_configure[21][12] ), .A2(n1196), .B1(
        \gpio_configure[27][12] ), .B2(n1198), .ZN(n909) );
  nr02d1 U1537 ( .A1(n905), .A2(n901), .ZN(n1166) );
  nr02d1 U1538 ( .A1(n900), .A2(n899), .ZN(n1191) );
  aoi22d1 U1539 ( .A1(\gpio_configure[17][12] ), .A2(n1166), .B1(
        \gpio_configure[10][12] ), .B2(n1191), .ZN(n908) );
  nr03d0 U1540 ( .A1(pad_count_1[4]), .A2(pad_count_1[3]), .A3(n1693), .ZN(
        n1146) );
  nr02d1 U1541 ( .A1(n903), .A2(n901), .ZN(n1199) );
  aoi22d1 U1542 ( .A1(\gpio_configure[0][12] ), .A2(n1146), .B1(
        \gpio_configure[19][12] ), .B2(n1199), .ZN(n907) );
  nr02d1 U1543 ( .A1(n903), .A2(n902), .ZN(n1175) );
  nr02d1 U1544 ( .A1(n905), .A2(n904), .ZN(n1174) );
  aoi22d1 U1545 ( .A1(\gpio_configure[31][12] ), .A2(n1175), .B1(
        \gpio_configure[5][12] ), .B2(n1174), .ZN(n906) );
  nr04d0 U1546 ( .A1(n913), .A2(n912), .A3(n911), .A4(n910), .ZN(n915) );
  inv0d0 U1547 ( .I(xfer_state[0]), .ZN(n1675) );
  nr02d0 U1548 ( .A1(n1675), .A2(xfer_state[1]), .ZN(n1696) );
  nd02d0 U1549 ( .A1(xfer_state[1]), .A2(n1675), .ZN(n1666) );
  nr02d1 U1550 ( .A1(n1649), .A2(n1666), .ZN(n1634) );
  inv0d1 U1551 ( .I(n1634), .ZN(n1476) );
  nd02d1 U1552 ( .A1(n1646), .A2(n1476), .ZN(n1214) );
  aoi22d1 U1553 ( .A1(serial_data_staging_1[12]), .A2(n1632), .B1(n1634), .B2(
        serial_data_staging_1[11]), .ZN(n914) );
  oai21d1 U1554 ( .B1(n915), .B2(n1646), .A(n914), .ZN(n2657) );
  nr02d0 U1555 ( .A1(xfer_count[3]), .A2(xfer_count[2]), .ZN(n1657) );
  inv0d0 U1556 ( .I(xfer_count[0]), .ZN(n1660) );
  nd02d0 U1557 ( .A1(xfer_state[1]), .A2(xfer_state[0]), .ZN(n1661) );
  aoi31d1 U1558 ( .B1(xfer_count[1]), .B2(n1657), .B3(n1660), .A(n1661), .ZN(
        n1658) );
  nd02d0 U1559 ( .A1(xfer_count[3]), .A2(xfer_count[2]), .ZN(n916) );
  nr03d0 U1560 ( .A1(xfer_count[0]), .A2(xfer_count[1]), .A3(n916), .ZN(n1651)
         );
  nd02d0 U1561 ( .A1(n1649), .A2(n1651), .ZN(n917) );
  or02d0 U1562 ( .A1(n1666), .A2(n917), .Z(n1645) );
  inv0d0 U1563 ( .I(xfer_state[1]), .ZN(n1687) );
  nd03d0 U1564 ( .A1(serial_xfer), .A2(n1687), .A3(n1675), .ZN(n1668) );
  nd13d1 U1565 ( .A1(n1658), .A2(n1645), .A3(n1668), .ZN(n2656) );
  inv0d0 U1566 ( .I(pad_count_2[1]), .ZN(n1672) );
  nr03d0 U1567 ( .A1(n1672), .A2(pad_count_2[4]), .A3(pad_count_2[3]), .ZN(
        n1216) );
  inv0d0 U1568 ( .I(pad_count_2[2]), .ZN(n1679) );
  inv0d0 U1569 ( .I(pad_count_2[5]), .ZN(n1683) );
  nr02d0 U1570 ( .A1(n1679), .A2(n1683), .ZN(n1559) );
  inv0d0 U1571 ( .I(pad_count_2[0]), .ZN(n1673) );
  aoi31d1 U1572 ( .B1(n1216), .B2(n1559), .B3(n1673), .A(n917), .ZN(n918) );
  nr02d0 U1573 ( .A1(n1696), .A2(n1658), .ZN(n1667) );
  oai21d1 U1574 ( .B1(n918), .B2(n1666), .A(n1667), .ZN(n2655) );
  aoi22d1 U1575 ( .A1(\gpio_configure[22][0] ), .A2(n1200), .B1(
        \gpio_configure[6][0] ), .B2(n1176), .ZN(n922) );
  aoi22d1 U1576 ( .A1(\gpio_configure[28][0] ), .A2(n1165), .B1(
        \gpio_configure[14][0] ), .B2(n1197), .ZN(n921) );
  aoi22d1 U1577 ( .A1(\gpio_configure[5][0] ), .A2(n1174), .B1(
        \gpio_configure[2][0] ), .B2(n1178), .ZN(n920) );
  aoi22d1 U1578 ( .A1(\gpio_configure[29][0] ), .A2(n1203), .B1(
        \gpio_configure[7][0] ), .B2(n1173), .ZN(n919) );
  aoi22d1 U1579 ( .A1(\gpio_configure[20][0] ), .A2(n1163), .B1(
        \gpio_configure[23][0] ), .B2(n1190), .ZN(n926) );
  aoi22d1 U1580 ( .A1(\gpio_configure[0][0] ), .A2(n1146), .B1(
        \gpio_configure[9][0] ), .B2(n1186), .ZN(n925) );
  aoi22d1 U1581 ( .A1(\gpio_configure[31][0] ), .A2(n1175), .B1(
        \gpio_configure[15][0] ), .B2(n1188), .ZN(n924) );
  aoi22d1 U1582 ( .A1(\gpio_configure[25][0] ), .A2(n1201), .B1(
        \gpio_configure[24][0] ), .B2(n1161), .ZN(n923) );
  aoi22d1 U1583 ( .A1(\gpio_configure[27][0] ), .A2(n1198), .B1(
        \gpio_configure[16][0] ), .B2(n1697), .ZN(n930) );
  aoi22d1 U1584 ( .A1(\gpio_configure[21][0] ), .A2(n1196), .B1(
        \gpio_configure[11][0] ), .B2(n1168), .ZN(n929) );
  aoi22d1 U1585 ( .A1(\gpio_configure[19][0] ), .A2(n1199), .B1(
        \gpio_configure[13][0] ), .B2(n1187), .ZN(n928) );
  aoi22d1 U1586 ( .A1(\gpio_configure[26][0] ), .A2(n1179), .B1(
        \gpio_configure[12][0] ), .B2(n1180), .ZN(n927) );
  aoi22d1 U1587 ( .A1(\gpio_configure[30][0] ), .A2(n1164), .B1(
        \gpio_configure[18][0] ), .B2(n1177), .ZN(n934) );
  aoi22d1 U1588 ( .A1(\gpio_configure[3][0] ), .A2(n1162), .B1(
        \gpio_configure[10][0] ), .B2(n1191), .ZN(n933) );
  aoi22d1 U1589 ( .A1(\gpio_configure[17][0] ), .A2(n1166), .B1(
        \gpio_configure[1][0] ), .B2(n1202), .ZN(n932) );
  aoi22d1 U1590 ( .A1(\gpio_configure[8][0] ), .A2(n1167), .B1(
        \gpio_configure[4][0] ), .B2(n1189), .ZN(n931) );
  nr04d0 U1591 ( .A1(n938), .A2(n937), .A3(n936), .A4(n935), .ZN(n939) );
  inv0d0 U1592 ( .I(serial_data_staging_1[0]), .ZN(n960) );
  oai22d1 U1593 ( .A1(n939), .A2(n1646), .B1(n1214), .B2(n960), .ZN(n2654) );
  inv0d0 U1594 ( .I(serial_data_staging_1[1]), .ZN(n982) );
  aoi22d1 U1595 ( .A1(\gpio_configure[31][1] ), .A2(n1175), .B1(
        \gpio_configure[13][1] ), .B2(n1187), .ZN(n943) );
  aoi22d1 U1596 ( .A1(\gpio_configure[4][1] ), .A2(n1189), .B1(
        \gpio_configure[2][1] ), .B2(n1178), .ZN(n942) );
  aoi22d1 U1597 ( .A1(\gpio_configure[30][1] ), .A2(n1164), .B1(
        \gpio_configure[29][1] ), .B2(n1203), .ZN(n941) );
  aoi22d1 U1598 ( .A1(\gpio_configure[23][1] ), .A2(n1190), .B1(
        \gpio_configure[11][1] ), .B2(n1168), .ZN(n940) );
  aoi22d1 U1599 ( .A1(\gpio_configure[28][1] ), .A2(n1165), .B1(
        \gpio_configure[6][1] ), .B2(n1176), .ZN(n947) );
  aoi22d1 U1600 ( .A1(\gpio_configure[18][1] ), .A2(n1177), .B1(
        \gpio_configure[25][1] ), .B2(n1201), .ZN(n946) );
  aoi22d1 U1601 ( .A1(\gpio_configure[21][1] ), .A2(n1196), .B1(
        \gpio_configure[5][1] ), .B2(n1174), .ZN(n945) );
  aoi22d1 U1602 ( .A1(\gpio_configure[20][1] ), .A2(n1163), .B1(
        \gpio_configure[22][1] ), .B2(n1200), .ZN(n944) );
  aoi22d1 U1603 ( .A1(\gpio_configure[3][1] ), .A2(n1162), .B1(
        \gpio_configure[14][1] ), .B2(n1197), .ZN(n951) );
  aoi22d1 U1604 ( .A1(\gpio_configure[16][1] ), .A2(n1697), .B1(
        \gpio_configure[7][1] ), .B2(n1173), .ZN(n950) );
  aoi22d1 U1605 ( .A1(\gpio_configure[0][1] ), .A2(n1146), .B1(
        \gpio_configure[9][1] ), .B2(n1186), .ZN(n949) );
  aoi22d1 U1606 ( .A1(\gpio_configure[19][1] ), .A2(n1199), .B1(
        \gpio_configure[12][1] ), .B2(n1180), .ZN(n948) );
  aoi22d1 U1607 ( .A1(\gpio_configure[17][1] ), .A2(n1166), .B1(
        \gpio_configure[10][1] ), .B2(n1191), .ZN(n955) );
  aoi22d1 U1608 ( .A1(\gpio_configure[24][1] ), .A2(n1161), .B1(
        \gpio_configure[26][1] ), .B2(n1179), .ZN(n954) );
  aoi22d1 U1609 ( .A1(\gpio_configure[15][1] ), .A2(n1188), .B1(
        \gpio_configure[1][1] ), .B2(n1202), .ZN(n953) );
  aoi22d1 U1610 ( .A1(\gpio_configure[27][1] ), .A2(n1198), .B1(
        \gpio_configure[8][1] ), .B2(n1167), .ZN(n952) );
  oai222d1 U1611 ( .A1(n982), .A2(n1214), .B1(n1646), .B2(n961), .C1(n1476), 
        .C2(n960), .ZN(n2653) );
  inv0d0 U1612 ( .I(serial_data_staging_1[2]), .ZN(n1004) );
  aoi22d1 U1613 ( .A1(\gpio_configure[9][2] ), .A2(n1186), .B1(
        \gpio_configure[11][2] ), .B2(n1168), .ZN(n965) );
  aoi22d1 U1614 ( .A1(\gpio_configure[29][2] ), .A2(n1203), .B1(
        \gpio_configure[2][2] ), .B2(n1178), .ZN(n964) );
  aoi22d1 U1615 ( .A1(\gpio_configure[24][2] ), .A2(n1161), .B1(
        \gpio_configure[8][2] ), .B2(n1167), .ZN(n963) );
  aoi22d1 U1616 ( .A1(\gpio_configure[23][2] ), .A2(n1190), .B1(
        \gpio_configure[5][2] ), .B2(n1174), .ZN(n962) );
  aoi22d1 U1617 ( .A1(\gpio_configure[6][2] ), .A2(n1176), .B1(
        \gpio_configure[3][2] ), .B2(n1162), .ZN(n969) );
  aoi22d1 U1618 ( .A1(\gpio_configure[27][2] ), .A2(n1198), .B1(
        \gpio_configure[20][2] ), .B2(n1163), .ZN(n968) );
  aoi22d1 U1619 ( .A1(\gpio_configure[0][2] ), .A2(n1146), .B1(
        \gpio_configure[4][2] ), .B2(n1189), .ZN(n967) );
  aoi22d1 U1620 ( .A1(\gpio_configure[21][2] ), .A2(n1196), .B1(
        \gpio_configure[1][2] ), .B2(n1202), .ZN(n966) );
  aoi22d1 U1621 ( .A1(\gpio_configure[19][2] ), .A2(n1199), .B1(
        \gpio_configure[7][2] ), .B2(n1173), .ZN(n973) );
  aoi22d1 U1622 ( .A1(\gpio_configure[30][2] ), .A2(n1164), .B1(
        \gpio_configure[18][2] ), .B2(n1177), .ZN(n972) );
  aoi22d1 U1623 ( .A1(\gpio_configure[22][2] ), .A2(n1200), .B1(
        \gpio_configure[25][2] ), .B2(n1201), .ZN(n971) );
  aoi22d1 U1624 ( .A1(\gpio_configure[28][2] ), .A2(n1165), .B1(
        \gpio_configure[16][2] ), .B2(n1697), .ZN(n970) );
  aoi22d1 U1625 ( .A1(\gpio_configure[31][2] ), .A2(n1175), .B1(
        \gpio_configure[17][2] ), .B2(n1166), .ZN(n977) );
  aoi22d1 U1626 ( .A1(\gpio_configure[10][2] ), .A2(n1191), .B1(
        \gpio_configure[12][2] ), .B2(n1180), .ZN(n976) );
  aoi22d1 U1627 ( .A1(\gpio_configure[14][2] ), .A2(n1197), .B1(
        \gpio_configure[15][2] ), .B2(n1188), .ZN(n975) );
  aoi22d1 U1628 ( .A1(\gpio_configure[26][2] ), .A2(n1179), .B1(
        \gpio_configure[13][2] ), .B2(n1187), .ZN(n974) );
  nr04d0 U1629 ( .A1(n981), .A2(n980), .A3(n979), .A4(n978), .ZN(n983) );
  oai222d1 U1630 ( .A1(n1004), .A2(n1214), .B1(n1646), .B2(n983), .C1(n1476), 
        .C2(n982), .ZN(n2652) );
  inv0d0 U1631 ( .I(serial_data_staging_1[3]), .ZN(n1026) );
  aoi22d1 U1632 ( .A1(\gpio_configure[27][3] ), .A2(n1198), .B1(
        \gpio_configure[21][3] ), .B2(n1196), .ZN(n987) );
  aoi22d1 U1633 ( .A1(\gpio_configure[20][3] ), .A2(n1163), .B1(
        \gpio_configure[14][3] ), .B2(n1197), .ZN(n986) );
  aoi22d1 U1634 ( .A1(\gpio_configure[18][3] ), .A2(n1177), .B1(
        \gpio_configure[6][3] ), .B2(n1176), .ZN(n985) );
  aoi22d1 U1635 ( .A1(\gpio_configure[19][3] ), .A2(n1199), .B1(
        \gpio_configure[3][3] ), .B2(n1162), .ZN(n984) );
  aoi22d1 U1636 ( .A1(\gpio_configure[9][3] ), .A2(n1186), .B1(
        \gpio_configure[16][3] ), .B2(n1697), .ZN(n991) );
  aoi22d1 U1637 ( .A1(\gpio_configure[28][3] ), .A2(n1165), .B1(
        \gpio_configure[7][3] ), .B2(n1173), .ZN(n990) );
  aoi22d1 U1638 ( .A1(\gpio_configure[23][3] ), .A2(n1190), .B1(
        \gpio_configure[2][3] ), .B2(n1178), .ZN(n989) );
  aoi22d1 U1639 ( .A1(\gpio_configure[5][3] ), .A2(n1174), .B1(
        \gpio_configure[12][3] ), .B2(n1180), .ZN(n988) );
  buffd1 U1640 ( .I(n1146), .Z(n1185) );
  aoi22d1 U1641 ( .A1(\gpio_configure[31][3] ), .A2(n1175), .B1(
        \gpio_configure[0][3] ), .B2(n1185), .ZN(n995) );
  aoi22d1 U1642 ( .A1(\gpio_configure[17][3] ), .A2(n1166), .B1(
        \gpio_configure[24][3] ), .B2(n1161), .ZN(n994) );
  aoi22d1 U1643 ( .A1(\gpio_configure[30][3] ), .A2(n1164), .B1(
        \gpio_configure[10][3] ), .B2(n1191), .ZN(n993) );
  aoi22d1 U1644 ( .A1(\gpio_configure[29][3] ), .A2(n1203), .B1(
        \gpio_configure[11][3] ), .B2(n1168), .ZN(n992) );
  aoi22d1 U1645 ( .A1(\gpio_configure[8][3] ), .A2(n1167), .B1(
        \gpio_configure[13][3] ), .B2(n1187), .ZN(n999) );
  aoi22d1 U1646 ( .A1(\gpio_configure[26][3] ), .A2(n1179), .B1(
        \gpio_configure[4][3] ), .B2(n1189), .ZN(n998) );
  aoi22d1 U1647 ( .A1(\gpio_configure[22][3] ), .A2(n1200), .B1(
        \gpio_configure[15][3] ), .B2(n1188), .ZN(n997) );
  aoi22d1 U1648 ( .A1(\gpio_configure[25][3] ), .A2(n1201), .B1(
        \gpio_configure[1][3] ), .B2(n1202), .ZN(n996) );
  nr04d0 U1649 ( .A1(n1003), .A2(n1002), .A3(n1001), .A4(n1000), .ZN(n1005) );
  oai222d1 U1650 ( .A1(n1026), .A2(n1214), .B1(n1646), .B2(n1005), .C1(n1476), 
        .C2(n1004), .ZN(n2651) );
  inv0d0 U1651 ( .I(serial_data_staging_1[4]), .ZN(n1048) );
  aoi22d1 U1652 ( .A1(\gpio_configure[8][4] ), .A2(n1167), .B1(
        \gpio_configure[2][4] ), .B2(n1178), .ZN(n1009) );
  aoi22d1 U1653 ( .A1(\gpio_configure[27][4] ), .A2(n1198), .B1(
        \gpio_configure[14][4] ), .B2(n1197), .ZN(n1008) );
  aoi22d1 U1654 ( .A1(\gpio_configure[22][4] ), .A2(n1200), .B1(
        \gpio_configure[19][4] ), .B2(n1199), .ZN(n1007) );
  aoi22d1 U1655 ( .A1(\gpio_configure[24][4] ), .A2(n1161), .B1(
        \gpio_configure[4][4] ), .B2(n1189), .ZN(n1006) );
  aoi22d1 U1656 ( .A1(\gpio_configure[0][4] ), .A2(n1146), .B1(
        \gpio_configure[30][4] ), .B2(n1164), .ZN(n1013) );
  aoi22d1 U1657 ( .A1(\gpio_configure[5][4] ), .A2(n1174), .B1(
        \gpio_configure[15][4] ), .B2(n1188), .ZN(n1012) );
  aoi22d1 U1658 ( .A1(\gpio_configure[3][4] ), .A2(n1162), .B1(
        \gpio_configure[6][4] ), .B2(n1176), .ZN(n1011) );
  aoi22d1 U1659 ( .A1(\gpio_configure[25][4] ), .A2(n1201), .B1(
        \gpio_configure[1][4] ), .B2(n1202), .ZN(n1010) );
  aoi22d1 U1660 ( .A1(\gpio_configure[23][4] ), .A2(n1190), .B1(
        \gpio_configure[12][4] ), .B2(n1180), .ZN(n1017) );
  aoi22d1 U1661 ( .A1(\gpio_configure[26][4] ), .A2(n1179), .B1(
        \gpio_configure[16][4] ), .B2(n1697), .ZN(n1016) );
  aoi22d1 U1662 ( .A1(\gpio_configure[10][4] ), .A2(n1191), .B1(
        \gpio_configure[13][4] ), .B2(n1187), .ZN(n1015) );
  aoi22d1 U1663 ( .A1(\gpio_configure[20][4] ), .A2(n1163), .B1(
        \gpio_configure[7][4] ), .B2(n1173), .ZN(n1014) );
  aoi22d1 U1664 ( .A1(\gpio_configure[21][4] ), .A2(n1196), .B1(
        \gpio_configure[28][4] ), .B2(n1165), .ZN(n1021) );
  aoi22d1 U1665 ( .A1(\gpio_configure[31][4] ), .A2(n1175), .B1(
        \gpio_configure[18][4] ), .B2(n1177), .ZN(n1020) );
  aoi22d1 U1666 ( .A1(\gpio_configure[17][4] ), .A2(n1166), .B1(
        \gpio_configure[9][4] ), .B2(n1186), .ZN(n1019) );
  aoi22d1 U1667 ( .A1(\gpio_configure[29][4] ), .A2(n1203), .B1(
        \gpio_configure[11][4] ), .B2(n1168), .ZN(n1018) );
  nr04d0 U1668 ( .A1(n1025), .A2(n1024), .A3(n1023), .A4(n1022), .ZN(n1027) );
  oai222d1 U1669 ( .A1(n1048), .A2(n1214), .B1(n1646), .B2(n1027), .C1(n1476), 
        .C2(n1026), .ZN(n2650) );
  inv0d0 U1670 ( .I(serial_data_staging_1[5]), .ZN(n1070) );
  aoi22d1 U1671 ( .A1(\gpio_configure[2][5] ), .A2(n1178), .B1(
        \gpio_configure[30][5] ), .B2(n1164), .ZN(n1031) );
  aoi22d1 U1672 ( .A1(\gpio_configure[14][5] ), .A2(n1197), .B1(
        \gpio_configure[13][5] ), .B2(n1187), .ZN(n1030) );
  aoi22d1 U1673 ( .A1(\gpio_configure[5][5] ), .A2(n1174), .B1(
        \gpio_configure[16][5] ), .B2(n1697), .ZN(n1029) );
  aoi22d1 U1674 ( .A1(\gpio_configure[6][5] ), .A2(n1176), .B1(
        \gpio_configure[18][5] ), .B2(n1177), .ZN(n1028) );
  aoi22d1 U1675 ( .A1(\gpio_configure[28][5] ), .A2(n1165), .B1(
        \gpio_configure[0][5] ), .B2(n1185), .ZN(n1035) );
  aoi22d1 U1676 ( .A1(\gpio_configure[7][5] ), .A2(n1173), .B1(
        \gpio_configure[25][5] ), .B2(n1201), .ZN(n1034) );
  aoi22d1 U1677 ( .A1(\gpio_configure[27][5] ), .A2(n1198), .B1(
        \gpio_configure[19][5] ), .B2(n1199), .ZN(n1033) );
  aoi22d1 U1678 ( .A1(\gpio_configure[1][5] ), .A2(n1202), .B1(
        \gpio_configure[31][5] ), .B2(n1175), .ZN(n1032) );
  aoi22d1 U1679 ( .A1(\gpio_configure[9][5] ), .A2(n1186), .B1(
        \gpio_configure[21][5] ), .B2(n1196), .ZN(n1039) );
  aoi22d1 U1680 ( .A1(\gpio_configure[11][5] ), .A2(n1168), .B1(
        \gpio_configure[23][5] ), .B2(n1190), .ZN(n1038) );
  aoi22d1 U1681 ( .A1(\gpio_configure[29][5] ), .A2(n1203), .B1(
        \gpio_configure[24][5] ), .B2(n1161), .ZN(n1037) );
  aoi22d1 U1682 ( .A1(\gpio_configure[8][5] ), .A2(n1167), .B1(
        \gpio_configure[4][5] ), .B2(n1189), .ZN(n1036) );
  aoi22d1 U1683 ( .A1(\gpio_configure[12][5] ), .A2(n1180), .B1(
        \gpio_configure[15][5] ), .B2(n1188), .ZN(n1043) );
  aoi22d1 U1684 ( .A1(\gpio_configure[3][5] ), .A2(n1162), .B1(
        \gpio_configure[26][5] ), .B2(n1179), .ZN(n1042) );
  aoi22d1 U1685 ( .A1(\gpio_configure[22][5] ), .A2(n1200), .B1(
        \gpio_configure[17][5] ), .B2(n1166), .ZN(n1041) );
  aoi22d1 U1686 ( .A1(\gpio_configure[10][5] ), .A2(n1191), .B1(
        \gpio_configure[20][5] ), .B2(n1163), .ZN(n1040) );
  nr04d0 U1687 ( .A1(n1047), .A2(n1046), .A3(n1045), .A4(n1044), .ZN(n1049) );
  oai222d1 U1688 ( .A1(n1070), .A2(n1214), .B1(n1646), .B2(n1049), .C1(n1476), 
        .C2(n1048), .ZN(n2649) );
  inv0d0 U1689 ( .I(serial_data_staging_1[6]), .ZN(n1092) );
  aoi22d1 U1690 ( .A1(\gpio_configure[4][6] ), .A2(n1189), .B1(
        \gpio_configure[8][6] ), .B2(n1167), .ZN(n1053) );
  aoi22d1 U1691 ( .A1(\gpio_configure[7][6] ), .A2(n1173), .B1(
        \gpio_configure[26][6] ), .B2(n1179), .ZN(n1052) );
  aoi22d1 U1692 ( .A1(\gpio_configure[9][6] ), .A2(n1186), .B1(
        \gpio_configure[18][6] ), .B2(n1177), .ZN(n1051) );
  aoi22d1 U1693 ( .A1(\gpio_configure[16][6] ), .A2(n1697), .B1(
        \gpio_configure[24][6] ), .B2(n1161), .ZN(n1050) );
  aoi22d1 U1694 ( .A1(\gpio_configure[13][6] ), .A2(n1187), .B1(
        \gpio_configure[2][6] ), .B2(n1178), .ZN(n1057) );
  aoi22d1 U1695 ( .A1(\gpio_configure[3][6] ), .A2(n1162), .B1(
        \gpio_configure[30][6] ), .B2(n1164), .ZN(n1056) );
  aoi22d1 U1696 ( .A1(\gpio_configure[12][6] ), .A2(n1180), .B1(
        \gpio_configure[1][6] ), .B2(n1202), .ZN(n1055) );
  aoi22d1 U1697 ( .A1(\gpio_configure[27][6] ), .A2(n1198), .B1(
        \gpio_configure[19][6] ), .B2(n1199), .ZN(n1054) );
  aoi22d1 U1698 ( .A1(\gpio_configure[11][6] ), .A2(n1168), .B1(
        \gpio_configure[31][6] ), .B2(n1175), .ZN(n1061) );
  aoi22d1 U1699 ( .A1(\gpio_configure[6][6] ), .A2(n1176), .B1(
        \gpio_configure[28][6] ), .B2(n1165), .ZN(n1060) );
  aoi22d1 U1700 ( .A1(\gpio_configure[25][6] ), .A2(n1201), .B1(
        \gpio_configure[23][6] ), .B2(n1190), .ZN(n1059) );
  aoi22d1 U1701 ( .A1(\gpio_configure[15][6] ), .A2(n1188), .B1(
        \gpio_configure[0][6] ), .B2(n1185), .ZN(n1058) );
  aoi22d1 U1702 ( .A1(\gpio_configure[14][6] ), .A2(n1197), .B1(
        \gpio_configure[29][6] ), .B2(n1203), .ZN(n1065) );
  aoi22d1 U1703 ( .A1(\gpio_configure[5][6] ), .A2(n1174), .B1(
        \gpio_configure[17][6] ), .B2(n1166), .ZN(n1064) );
  aoi22d1 U1704 ( .A1(\gpio_configure[21][6] ), .A2(n1196), .B1(
        \gpio_configure[22][6] ), .B2(n1200), .ZN(n1063) );
  aoi22d1 U1705 ( .A1(\gpio_configure[10][6] ), .A2(n1191), .B1(
        \gpio_configure[20][6] ), .B2(n1163), .ZN(n1062) );
  nr04d0 U1706 ( .A1(n1069), .A2(n1068), .A3(n1067), .A4(n1066), .ZN(n1071) );
  oai222d1 U1707 ( .A1(n1092), .A2(n1214), .B1(n1646), .B2(n1071), .C1(n1476), 
        .C2(n1070), .ZN(n2648) );
  inv0d0 U1708 ( .I(serial_data_staging_1[7]), .ZN(n1114) );
  aoi22d1 U1709 ( .A1(\gpio_configure[14][7] ), .A2(n1197), .B1(
        \gpio_configure[24][7] ), .B2(n1161), .ZN(n1075) );
  aoi22d1 U1710 ( .A1(\gpio_configure[10][7] ), .A2(n1191), .B1(
        \gpio_configure[22][7] ), .B2(n1200), .ZN(n1074) );
  aoi22d1 U1711 ( .A1(\gpio_configure[9][7] ), .A2(n1186), .B1(
        \gpio_configure[3][7] ), .B2(n1162), .ZN(n1073) );
  aoi22d1 U1712 ( .A1(\gpio_configure[13][7] ), .A2(n1187), .B1(
        \gpio_configure[17][7] ), .B2(n1166), .ZN(n1072) );
  aoi22d1 U1713 ( .A1(\gpio_configure[26][7] ), .A2(n1179), .B1(
        \gpio_configure[30][7] ), .B2(n1164), .ZN(n1079) );
  aoi22d1 U1714 ( .A1(\gpio_configure[8][7] ), .A2(n1167), .B1(
        \gpio_configure[15][7] ), .B2(n1188), .ZN(n1078) );
  aoi22d1 U1715 ( .A1(\gpio_configure[6][7] ), .A2(n1176), .B1(
        \gpio_configure[18][7] ), .B2(n1177), .ZN(n1077) );
  aoi22d1 U1716 ( .A1(\gpio_configure[7][7] ), .A2(n1173), .B1(
        \gpio_configure[0][7] ), .B2(n1185), .ZN(n1076) );
  aoi22d1 U1717 ( .A1(\gpio_configure[23][7] ), .A2(n1190), .B1(
        \gpio_configure[29][7] ), .B2(n1203), .ZN(n1083) );
  aoi22d1 U1718 ( .A1(\gpio_configure[11][7] ), .A2(n1168), .B1(
        \gpio_configure[5][7] ), .B2(n1174), .ZN(n1082) );
  aoi22d1 U1719 ( .A1(\gpio_configure[4][7] ), .A2(n1189), .B1(
        \gpio_configure[21][7] ), .B2(n1196), .ZN(n1081) );
  aoi22d1 U1720 ( .A1(\gpio_configure[27][7] ), .A2(n1198), .B1(
        \gpio_configure[28][7] ), .B2(n1165), .ZN(n1080) );
  aoi22d1 U1721 ( .A1(\gpio_configure[1][7] ), .A2(n1202), .B1(
        \gpio_configure[16][7] ), .B2(n1697), .ZN(n1087) );
  aoi22d1 U1722 ( .A1(\gpio_configure[2][7] ), .A2(n1178), .B1(
        \gpio_configure[31][7] ), .B2(n1175), .ZN(n1086) );
  aoi22d1 U1723 ( .A1(\gpio_configure[12][7] ), .A2(n1180), .B1(
        \gpio_configure[20][7] ), .B2(n1163), .ZN(n1085) );
  aoi22d1 U1724 ( .A1(\gpio_configure[19][7] ), .A2(n1199), .B1(
        \gpio_configure[25][7] ), .B2(n1201), .ZN(n1084) );
  nr04d0 U1725 ( .A1(n1091), .A2(n1090), .A3(n1089), .A4(n1088), .ZN(n1093) );
  oai222d1 U1726 ( .A1(n1114), .A2(n1214), .B1(n1646), .B2(n1093), .C1(n1476), 
        .C2(n1092), .ZN(n2647) );
  inv0d0 U1727 ( .I(serial_data_staging_1[8]), .ZN(n1136) );
  aoi22d1 U1728 ( .A1(\gpio_configure[29][8] ), .A2(n1203), .B1(
        \gpio_configure[16][8] ), .B2(n1697), .ZN(n1097) );
  aoi22d1 U1729 ( .A1(\gpio_configure[20][8] ), .A2(n1163), .B1(
        \gpio_configure[2][8] ), .B2(n1178), .ZN(n1096) );
  aoi22d1 U1730 ( .A1(\gpio_configure[21][8] ), .A2(n1196), .B1(
        \gpio_configure[1][8] ), .B2(n1202), .ZN(n1095) );
  aoi22d1 U1731 ( .A1(\gpio_configure[26][8] ), .A2(n1179), .B1(
        \gpio_configure[11][8] ), .B2(n1168), .ZN(n1094) );
  aoi22d1 U1732 ( .A1(\gpio_configure[5][8] ), .A2(n1174), .B1(
        \gpio_configure[10][8] ), .B2(n1191), .ZN(n1101) );
  aoi22d1 U1733 ( .A1(\gpio_configure[30][8] ), .A2(n1164), .B1(
        \gpio_configure[7][8] ), .B2(n1173), .ZN(n1100) );
  aoi22d1 U1734 ( .A1(\gpio_configure[24][8] ), .A2(n1161), .B1(
        \gpio_configure[14][8] ), .B2(n1197), .ZN(n1099) );
  aoi22d1 U1735 ( .A1(\gpio_configure[23][8] ), .A2(n1190), .B1(
        \gpio_configure[17][8] ), .B2(n1166), .ZN(n1098) );
  aoi22d1 U1736 ( .A1(\gpio_configure[28][8] ), .A2(n1165), .B1(
        \gpio_configure[3][8] ), .B2(n1162), .ZN(n1105) );
  aoi22d1 U1737 ( .A1(\gpio_configure[25][8] ), .A2(n1201), .B1(
        \gpio_configure[0][8] ), .B2(n1185), .ZN(n1104) );
  aoi22d1 U1738 ( .A1(\gpio_configure[27][8] ), .A2(n1198), .B1(
        \gpio_configure[31][8] ), .B2(n1175), .ZN(n1103) );
  aoi22d1 U1739 ( .A1(\gpio_configure[4][8] ), .A2(n1189), .B1(
        \gpio_configure[8][8] ), .B2(n1167), .ZN(n1102) );
  aoi22d1 U1740 ( .A1(\gpio_configure[22][8] ), .A2(n1200), .B1(
        \gpio_configure[15][8] ), .B2(n1188), .ZN(n1109) );
  aoi22d1 U1741 ( .A1(\gpio_configure[18][8] ), .A2(n1177), .B1(
        \gpio_configure[6][8] ), .B2(n1176), .ZN(n1108) );
  aoi22d1 U1742 ( .A1(\gpio_configure[12][8] ), .A2(n1180), .B1(
        \gpio_configure[9][8] ), .B2(n1186), .ZN(n1107) );
  aoi22d1 U1743 ( .A1(\gpio_configure[19][8] ), .A2(n1199), .B1(
        \gpio_configure[13][8] ), .B2(n1187), .ZN(n1106) );
  oai222d1 U1744 ( .A1(n1136), .A2(n1214), .B1(n1646), .B2(n1115), .C1(n1476), 
        .C2(n1114), .ZN(n2646) );
  inv0d0 U1745 ( .I(serial_data_staging_1[9]), .ZN(n1159) );
  aoi22d1 U1746 ( .A1(\gpio_configure[5][9] ), .A2(n1174), .B1(
        \gpio_configure[21][9] ), .B2(n1196), .ZN(n1119) );
  aoi22d1 U1747 ( .A1(\gpio_configure[9][9] ), .A2(n1186), .B1(
        \gpio_configure[31][9] ), .B2(n1175), .ZN(n1118) );
  aoi22d1 U1748 ( .A1(\gpio_configure[16][9] ), .A2(n1697), .B1(
        \gpio_configure[8][9] ), .B2(n1167), .ZN(n1117) );
  aoi22d1 U1749 ( .A1(\gpio_configure[28][9] ), .A2(n1165), .B1(
        \gpio_configure[27][9] ), .B2(n1198), .ZN(n1116) );
  aoi22d1 U1750 ( .A1(\gpio_configure[4][9] ), .A2(n1189), .B1(
        \gpio_configure[30][9] ), .B2(n1164), .ZN(n1123) );
  aoi22d1 U1751 ( .A1(\gpio_configure[22][9] ), .A2(n1200), .B1(
        \gpio_configure[20][9] ), .B2(n1163), .ZN(n1122) );
  aoi22d1 U1752 ( .A1(\gpio_configure[2][9] ), .A2(n1178), .B1(
        \gpio_configure[11][9] ), .B2(n1168), .ZN(n1121) );
  aoi22d1 U1753 ( .A1(\gpio_configure[3][9] ), .A2(n1162), .B1(
        \gpio_configure[1][9] ), .B2(n1202), .ZN(n1120) );
  aoi22d1 U1754 ( .A1(\gpio_configure[6][9] ), .A2(n1176), .B1(
        \gpio_configure[29][9] ), .B2(n1203), .ZN(n1127) );
  aoi22d1 U1755 ( .A1(\gpio_configure[7][9] ), .A2(n1173), .B1(
        \gpio_configure[18][9] ), .B2(n1177), .ZN(n1126) );
  aoi22d1 U1756 ( .A1(\gpio_configure[12][9] ), .A2(n1180), .B1(
        \gpio_configure[13][9] ), .B2(n1187), .ZN(n1125) );
  aoi22d1 U1757 ( .A1(\gpio_configure[14][9] ), .A2(n1197), .B1(
        \gpio_configure[15][9] ), .B2(n1188), .ZN(n1124) );
  aoi22d1 U1758 ( .A1(\gpio_configure[23][9] ), .A2(n1190), .B1(
        \gpio_configure[0][9] ), .B2(n1185), .ZN(n1131) );
  aoi22d1 U1759 ( .A1(\gpio_configure[17][9] ), .A2(n1166), .B1(
        \gpio_configure[19][9] ), .B2(n1199), .ZN(n1130) );
  aoi22d1 U1760 ( .A1(\gpio_configure[10][9] ), .A2(n1191), .B1(
        \gpio_configure[25][9] ), .B2(n1201), .ZN(n1129) );
  aoi22d1 U1761 ( .A1(\gpio_configure[26][9] ), .A2(n1179), .B1(
        \gpio_configure[24][9] ), .B2(n1161), .ZN(n1128) );
  nr04d0 U1762 ( .A1(n1135), .A2(n1134), .A3(n1133), .A4(n1132), .ZN(n1137) );
  oai222d1 U1763 ( .A1(n1159), .A2(n1214), .B1(n1646), .B2(n1137), .C1(n1476), 
        .C2(n1136), .ZN(n2645) );
  inv0d0 U1764 ( .I(serial_data_staging_1[10]), .ZN(n1212) );
  aoi22d1 U1765 ( .A1(\gpio_configure[25][10] ), .A2(n1201), .B1(
        \gpio_configure[28][10] ), .B2(n1165), .ZN(n1141) );
  aoi22d1 U1766 ( .A1(\gpio_configure[26][10] ), .A2(n1179), .B1(
        \gpio_configure[8][10] ), .B2(n1167), .ZN(n1140) );
  aoi22d1 U1767 ( .A1(\gpio_configure[22][10] ), .A2(n1200), .B1(
        \gpio_configure[9][10] ), .B2(n1186), .ZN(n1139) );
  aoi22d1 U1768 ( .A1(\gpio_configure[27][10] ), .A2(n1198), .B1(
        \gpio_configure[3][10] ), .B2(n1162), .ZN(n1138) );
  aoi22d1 U1769 ( .A1(\gpio_configure[21][10] ), .A2(n1196), .B1(
        \gpio_configure[13][10] ), .B2(n1187), .ZN(n1145) );
  aoi22d1 U1770 ( .A1(\gpio_configure[30][10] ), .A2(n1164), .B1(
        \gpio_configure[17][10] ), .B2(n1166), .ZN(n1144) );
  aoi22d1 U1771 ( .A1(\gpio_configure[19][10] ), .A2(n1199), .B1(
        \gpio_configure[15][10] ), .B2(n1188), .ZN(n1143) );
  aoi22d1 U1772 ( .A1(\gpio_configure[23][10] ), .A2(n1190), .B1(
        \gpio_configure[4][10] ), .B2(n1189), .ZN(n1142) );
  aoi22d1 U1773 ( .A1(\gpio_configure[14][10] ), .A2(n1197), .B1(
        \gpio_configure[11][10] ), .B2(n1168), .ZN(n1150) );
  aoi22d1 U1774 ( .A1(\gpio_configure[24][10] ), .A2(n1161), .B1(
        \gpio_configure[7][10] ), .B2(n1173), .ZN(n1149) );
  aoi22d1 U1775 ( .A1(\gpio_configure[0][10] ), .A2(n1146), .B1(
        \gpio_configure[2][10] ), .B2(n1178), .ZN(n1148) );
  aoi22d1 U1776 ( .A1(\gpio_configure[1][10] ), .A2(n1202), .B1(
        \gpio_configure[10][10] ), .B2(n1191), .ZN(n1147) );
  aoi22d1 U1777 ( .A1(\gpio_configure[29][10] ), .A2(n1203), .B1(
        \gpio_configure[5][10] ), .B2(n1174), .ZN(n1154) );
  aoi22d1 U1778 ( .A1(\gpio_configure[6][10] ), .A2(n1176), .B1(
        \gpio_configure[16][10] ), .B2(n1697), .ZN(n1153) );
  aoi22d1 U1779 ( .A1(\gpio_configure[20][10] ), .A2(n1163), .B1(
        \gpio_configure[12][10] ), .B2(n1180), .ZN(n1152) );
  aoi22d1 U1780 ( .A1(\gpio_configure[18][10] ), .A2(n1177), .B1(
        \gpio_configure[31][10] ), .B2(n1175), .ZN(n1151) );
  nr04d0 U1781 ( .A1(n1158), .A2(n1157), .A3(n1156), .A4(n1155), .ZN(n1160) );
  oai222d1 U1782 ( .A1(n1212), .A2(n1214), .B1(n1646), .B2(n1160), .C1(n1476), 
        .C2(n1159), .ZN(n2644) );
  inv0d0 U1783 ( .I(serial_data_staging_1[11]), .ZN(n1215) );
  aoi22d1 U1784 ( .A1(\gpio_configure[3][11] ), .A2(n1162), .B1(
        \gpio_configure[24][11] ), .B2(n1161), .ZN(n1172) );
  aoi22d1 U1785 ( .A1(\gpio_configure[30][11] ), .A2(n1164), .B1(
        \gpio_configure[20][11] ), .B2(n1163), .ZN(n1171) );
  aoi22d1 U1786 ( .A1(\gpio_configure[17][11] ), .A2(n1166), .B1(
        \gpio_configure[28][11] ), .B2(n1165), .ZN(n1170) );
  aoi22d1 U1787 ( .A1(\gpio_configure[11][11] ), .A2(n1168), .B1(
        \gpio_configure[8][11] ), .B2(n1167), .ZN(n1169) );
  aoi22d1 U1788 ( .A1(\gpio_configure[5][11] ), .A2(n1174), .B1(
        \gpio_configure[7][11] ), .B2(n1173), .ZN(n1184) );
  aoi22d1 U1789 ( .A1(\gpio_configure[6][11] ), .A2(n1176), .B1(
        \gpio_configure[31][11] ), .B2(n1175), .ZN(n1183) );
  aoi22d1 U1790 ( .A1(\gpio_configure[2][11] ), .A2(n1178), .B1(
        \gpio_configure[18][11] ), .B2(n1177), .ZN(n1182) );
  aoi22d1 U1791 ( .A1(\gpio_configure[12][11] ), .A2(n1180), .B1(
        \gpio_configure[26][11] ), .B2(n1179), .ZN(n1181) );
  aoi22d1 U1792 ( .A1(\gpio_configure[9][11] ), .A2(n1186), .B1(
        \gpio_configure[0][11] ), .B2(n1185), .ZN(n1195) );
  aoi22d1 U1793 ( .A1(\gpio_configure[15][11] ), .A2(n1188), .B1(
        \gpio_configure[13][11] ), .B2(n1187), .ZN(n1194) );
  aoi22d1 U1794 ( .A1(\gpio_configure[16][11] ), .A2(n1697), .B1(
        \gpio_configure[4][11] ), .B2(n1189), .ZN(n1193) );
  aoi22d1 U1795 ( .A1(\gpio_configure[10][11] ), .A2(n1191), .B1(
        \gpio_configure[23][11] ), .B2(n1190), .ZN(n1192) );
  aoi22d1 U1796 ( .A1(\gpio_configure[14][11] ), .A2(n1197), .B1(
        \gpio_configure[21][11] ), .B2(n1196), .ZN(n1207) );
  aoi22d1 U1797 ( .A1(\gpio_configure[19][11] ), .A2(n1199), .B1(
        \gpio_configure[27][11] ), .B2(n1198), .ZN(n1206) );
  aoi22d1 U1798 ( .A1(\gpio_configure[25][11] ), .A2(n1201), .B1(
        \gpio_configure[22][11] ), .B2(n1200), .ZN(n1205) );
  aoi22d1 U1799 ( .A1(\gpio_configure[29][11] ), .A2(n1203), .B1(
        \gpio_configure[1][11] ), .B2(n1202), .ZN(n1204) );
  nr04d0 U1800 ( .A1(n1211), .A2(n1210), .A3(n1209), .A4(n1208), .ZN(n1213) );
  oai222d1 U1801 ( .A1(n1215), .A2(n1214), .B1(n1646), .B2(n1213), .C1(n1476), 
        .C2(n1212), .ZN(n2643) );
  nd03d0 U1802 ( .A1(pad_count_2[0]), .A2(n1679), .A3(n1683), .ZN(n1236) );
  nd03d0 U1803 ( .A1(pad_count_2[4]), .A2(pad_count_2[3]), .A3(pad_count_2[1]), 
        .ZN(n1678) );
  nr02d1 U1804 ( .A1(n1236), .A2(n1678), .ZN(n1591) );
  nd03d0 U1805 ( .A1(pad_count_2[2]), .A2(n1673), .A3(n1683), .ZN(n1234) );
  inv0d0 U1806 ( .I(pad_count_2[4]), .ZN(n1682) );
  nd03d0 U1807 ( .A1(pad_count_2[3]), .A2(n1682), .A3(n1672), .ZN(n1235) );
  nr02d1 U1808 ( .A1(n1234), .A2(n1235), .ZN(n1612) );
  aoi22d1 U1809 ( .A1(\gpio_configure[27][0] ), .A2(n1591), .B1(
        \gpio_configure[12][0] ), .B2(n1612), .ZN(n1220) );
  nd03d0 U1810 ( .A1(pad_count_2[3]), .A2(pad_count_2[1]), .A3(n1682), .ZN(
        n1239) );
  nr02d1 U1811 ( .A1(n1239), .A2(n1236), .ZN(n1607) );
  inv0d0 U1812 ( .I(n1216), .ZN(n1226) );
  nr02d1 U1813 ( .A1(n1231), .A2(n1226), .ZN(n1583) );
  aoi22d1 U1814 ( .A1(\gpio_configure[11][0] ), .A2(n1607), .B1(
        \gpio_configure[2][0] ), .B2(n1583), .ZN(n1219) );
  inv0d0 U1815 ( .I(pad_count_2[3]), .ZN(n1676) );
  nd03d0 U1816 ( .A1(pad_count_2[4]), .A2(pad_count_2[1]), .A3(n1676), .ZN(
        n1232) );
  nd03d0 U1817 ( .A1(pad_count_2[0]), .A2(pad_count_2[2]), .A3(n1683), .ZN(
        n1238) );
  nr02d1 U1818 ( .A1(n1232), .A2(n1238), .ZN(n1615) );
  nd03d0 U1819 ( .A1(pad_count_2[3]), .A2(pad_count_2[4]), .A3(n1672), .ZN(
        n1237) );
  nr02d1 U1820 ( .A1(n1237), .A2(n1234), .ZN(n1604) );
  aoi22d1 U1821 ( .A1(\gpio_configure[23][0] ), .A2(n1615), .B1(
        \gpio_configure[28][0] ), .B2(n1604), .ZN(n1218) );
  nr02d1 U1822 ( .A1(n1232), .A2(n1236), .ZN(n1577) );
  nr02d1 U1823 ( .A1(n1238), .A2(n1225), .ZN(n1618) );
  aoi22d1 U1824 ( .A1(\gpio_configure[19][0] ), .A2(n1577), .B1(
        \gpio_configure[5][0] ), .B2(n1618), .ZN(n1217) );
  nr02d1 U1825 ( .A1(n1237), .A2(n1238), .ZN(n1617) );
  nr02d1 U1826 ( .A1(n1231), .A2(n1239), .ZN(n1616) );
  aoi22d1 U1827 ( .A1(\gpio_configure[29][0] ), .A2(n1617), .B1(
        \gpio_configure[10][0] ), .B2(n1616), .ZN(n1224) );
  nr02d1 U1828 ( .A1(n1238), .A2(n1226), .ZN(n1600) );
  nr02d1 U1829 ( .A1(n1235), .A2(n1238), .ZN(n1582) );
  aoi22d1 U1830 ( .A1(\gpio_configure[7][0] ), .A2(n1600), .B1(
        \gpio_configure[13][0] ), .B2(n1582), .ZN(n1223) );
  nr02d1 U1831 ( .A1(n1234), .A2(n1226), .ZN(n1602) );
  nr02d1 U1832 ( .A1(n1231), .A2(n1235), .ZN(n1578) );
  aoi22d1 U1833 ( .A1(\gpio_configure[6][0] ), .A2(n1602), .B1(
        \gpio_configure[8][0] ), .B2(n1578), .ZN(n1222) );
  nr02d1 U1834 ( .A1(n1238), .A2(n1678), .ZN(n1601) );
  nd03d0 U1835 ( .A1(pad_count_2[4]), .A2(n1676), .A3(n1672), .ZN(n1233) );
  nr02d1 U1836 ( .A1(n1231), .A2(n1233), .ZN(n1606) );
  aoi22d1 U1837 ( .A1(\gpio_configure[31][0] ), .A2(n1601), .B1(
        \gpio_configure[16][0] ), .B2(n1606), .ZN(n1221) );
  nr02d1 U1838 ( .A1(n1234), .A2(n1239), .ZN(n1594) );
  nr02d1 U1839 ( .A1(n1236), .A2(n1225), .ZN(n1605) );
  aoi22d1 U1840 ( .A1(\gpio_configure[14][0] ), .A2(n1594), .B1(
        \gpio_configure[1][0] ), .B2(n1605), .ZN(n1230) );
  nr02d1 U1841 ( .A1(n1231), .A2(n1237), .ZN(n1579) );
  nr02d1 U1842 ( .A1(n1234), .A2(n1225), .ZN(n1590) );
  aoi22d1 U1843 ( .A1(\gpio_configure[24][0] ), .A2(n1579), .B1(
        \gpio_configure[4][0] ), .B2(n1590), .ZN(n1229) );
  nr02d1 U1844 ( .A1(n1234), .A2(n1678), .ZN(n1619) );
  nr02d1 U1845 ( .A1(n1238), .A2(n1233), .ZN(n1593) );
  aoi22d1 U1846 ( .A1(\gpio_configure[30][0] ), .A2(n1619), .B1(
        \gpio_configure[21][0] ), .B2(n1593), .ZN(n1228) );
  nr02d1 U1847 ( .A1(n1231), .A2(n1225), .ZN(n1581) );
  nr02d1 U1848 ( .A1(n1236), .A2(n1226), .ZN(n1613) );
  aoi22d1 U1849 ( .A1(\gpio_configure[0][0] ), .A2(n1581), .B1(
        \gpio_configure[3][0] ), .B2(n1613), .ZN(n1227) );
  nr02d1 U1850 ( .A1(n1231), .A2(n1678), .ZN(n1592) );
  nr02d1 U1851 ( .A1(n1231), .A2(n1232), .ZN(n1580) );
  aoi22d1 U1852 ( .A1(\gpio_configure[26][0] ), .A2(n1592), .B1(
        \gpio_configure[18][0] ), .B2(n1580), .ZN(n1243) );
  nr02d1 U1853 ( .A1(n1232), .A2(n1234), .ZN(n1589) );
  nr02d1 U1854 ( .A1(n1236), .A2(n1233), .ZN(n1576) );
  aoi22d1 U1855 ( .A1(\gpio_configure[22][0] ), .A2(n1589), .B1(
        \gpio_configure[17][0] ), .B2(n1576), .ZN(n1242) );
  nr02d1 U1856 ( .A1(n1234), .A2(n1233), .ZN(n1614) );
  nr02d1 U1857 ( .A1(n1236), .A2(n1235), .ZN(n1595) );
  aoi22d1 U1858 ( .A1(\gpio_configure[20][0] ), .A2(n1614), .B1(
        \gpio_configure[9][0] ), .B2(n1595), .ZN(n1241) );
  nr02d1 U1859 ( .A1(n1237), .A2(n1236), .ZN(n1603) );
  nr02d1 U1860 ( .A1(n1239), .A2(n1238), .ZN(n1588) );
  aoi22d1 U1861 ( .A1(\gpio_configure[25][0] ), .A2(n1603), .B1(
        \gpio_configure[15][0] ), .B2(n1588), .ZN(n1240) );
  nr04d0 U1862 ( .A1(n1247), .A2(n1246), .A3(n1245), .A4(n1244), .ZN(n1255) );
  nr04d0 U1863 ( .A1(pad_count_2[0]), .A2(pad_count_2[2]), .A3(n1646), .A4(
        n1683), .ZN(n1446) );
  nd02d0 U1864 ( .A1(n1446), .A2(n1672), .ZN(n1638) );
  inv0d0 U1865 ( .I(n1638), .ZN(n1538) );
  aoi22d1 U1866 ( .A1(\gpio_configure[32][0] ), .A2(n1538), .B1(n1632), .B2(
        serial_data_staging_2[0]), .ZN(n1254) );
  inv0d0 U1867 ( .I(\gpio_configure[36][0] ), .ZN(n1252) );
  nd02d1 U1868 ( .A1(pad_count_2[1]), .A2(n1446), .ZN(n1628) );
  inv0d0 U1869 ( .I(n1628), .ZN(n1537) );
  nr02d0 U1870 ( .A1(n1646), .A2(n1673), .ZN(n1248) );
  nd04d0 U1871 ( .A1(n1679), .A2(n1672), .A3(pad_count_2[5]), .A4(n1248), .ZN(
        n1478) );
  inv0d0 U1872 ( .I(n1478), .ZN(n1633) );
  aoi22d1 U1873 ( .A1(\gpio_configure[34][0] ), .A2(n1537), .B1(
        \gpio_configure[33][0] ), .B2(n1633), .ZN(n1251) );
  inv0d0 U1874 ( .I(n1248), .ZN(n1670) );
  nr03d0 U1875 ( .A1(n1679), .A2(n1683), .A3(n1670), .ZN(n1635) );
  nd02d0 U1876 ( .A1(pad_count_2[1]), .A2(n1248), .ZN(n1677) );
  nr02d0 U1877 ( .A1(pad_count_2[2]), .A2(n1677), .ZN(n1249) );
  nd02d0 U1878 ( .A1(pad_count_2[5]), .A2(n1249), .ZN(n1630) );
  inv0d0 U1879 ( .I(n1630), .ZN(n1570) );
  aoi22d1 U1880 ( .A1(\gpio_configure[37][0] ), .A2(n1635), .B1(
        \gpio_configure[35][0] ), .B2(n1570), .ZN(n1250) );
  ora211d1 U1881 ( .C1(n1252), .C2(n1541), .A(n1251), .B(n1250), .Z(n1253) );
  oai211d1 U1882 ( .C1(n1255), .C2(n1646), .A(n1254), .B(n1253), .ZN(n2642) );
  aoi22d1 U1883 ( .A1(\gpio_configure[8][1] ), .A2(n1578), .B1(
        \gpio_configure[4][1] ), .B2(n1590), .ZN(n1259) );
  aoi22d1 U1884 ( .A1(\gpio_configure[27][1] ), .A2(n1591), .B1(
        \gpio_configure[15][1] ), .B2(n1588), .ZN(n1258) );
  aoi22d1 U1885 ( .A1(\gpio_configure[11][1] ), .A2(n1607), .B1(
        \gpio_configure[1][1] ), .B2(n1605), .ZN(n1257) );
  aoi22d1 U1886 ( .A1(\gpio_configure[12][1] ), .A2(n1612), .B1(
        \gpio_configure[2][1] ), .B2(n1583), .ZN(n1256) );
  aoi22d1 U1887 ( .A1(\gpio_configure[22][1] ), .A2(n1589), .B1(
        \gpio_configure[10][1] ), .B2(n1616), .ZN(n1263) );
  aoi22d1 U1888 ( .A1(\gpio_configure[30][1] ), .A2(n1619), .B1(
        \gpio_configure[7][1] ), .B2(n1600), .ZN(n1262) );
  aoi22d1 U1889 ( .A1(\gpio_configure[18][1] ), .A2(n1580), .B1(
        \gpio_configure[28][1] ), .B2(n1604), .ZN(n1261) );
  aoi22d1 U1890 ( .A1(\gpio_configure[16][1] ), .A2(n1606), .B1(
        \gpio_configure[9][1] ), .B2(n1595), .ZN(n1260) );
  aoi22d1 U1891 ( .A1(\gpio_configure[0][1] ), .A2(n1581), .B1(
        \gpio_configure[17][1] ), .B2(n1576), .ZN(n1267) );
  aoi22d1 U1892 ( .A1(\gpio_configure[19][1] ), .A2(n1577), .B1(
        \gpio_configure[3][1] ), .B2(n1613), .ZN(n1266) );
  aoi22d1 U1893 ( .A1(\gpio_configure[20][1] ), .A2(n1614), .B1(
        \gpio_configure[6][1] ), .B2(n1602), .ZN(n1265) );
  aoi22d1 U1894 ( .A1(\gpio_configure[23][1] ), .A2(n1615), .B1(
        \gpio_configure[31][1] ), .B2(n1601), .ZN(n1264) );
  aoi22d1 U1895 ( .A1(\gpio_configure[24][1] ), .A2(n1579), .B1(
        \gpio_configure[21][1] ), .B2(n1593), .ZN(n1271) );
  aoi22d1 U1896 ( .A1(\gpio_configure[26][1] ), .A2(n1592), .B1(
        \gpio_configure[5][1] ), .B2(n1618), .ZN(n1270) );
  aoi22d1 U1897 ( .A1(\gpio_configure[25][1] ), .A2(n1603), .B1(
        \gpio_configure[14][1] ), .B2(n1594), .ZN(n1269) );
  aoi22d1 U1898 ( .A1(\gpio_configure[29][1] ), .A2(n1617), .B1(
        \gpio_configure[13][1] ), .B2(n1582), .ZN(n1268) );
  nr04d0 U1899 ( .A1(n1275), .A2(n1274), .A3(n1273), .A4(n1272), .ZN(n1281) );
  aor22d1 U1900 ( .A1(\gpio_configure[35][1] ), .A2(n1570), .B1(
        \gpio_configure[37][1] ), .B2(n1635), .Z(n1279) );
  aoi22d1 U1901 ( .A1(\gpio_configure[32][1] ), .A2(n1538), .B1(n1632), .B2(
        serial_data_staging_2[1]), .ZN(n1277) );
  aoi22d1 U1902 ( .A1(\gpio_configure[36][1] ), .A2(n1642), .B1(n1634), .B2(
        serial_data_staging_2[0]), .ZN(n1276) );
  oaim211d1 U1903 ( .C1(\gpio_configure[34][1] ), .C2(n1537), .A(n1277), .B(
        n1276), .ZN(n1278) );
  aoi211d1 U1904 ( .C1(\gpio_configure[33][1] ), .C2(n1633), .A(n1279), .B(
        n1278), .ZN(n1280) );
  oai21d1 U1905 ( .B1(n1281), .B2(n1646), .A(n1280), .ZN(n2641) );
  aoi22d1 U1906 ( .A1(\gpio_configure[17][2] ), .A2(n1576), .B1(
        \gpio_configure[7][2] ), .B2(n1600), .ZN(n1285) );
  aoi22d1 U1907 ( .A1(\gpio_configure[29][2] ), .A2(n1617), .B1(
        \gpio_configure[15][2] ), .B2(n1588), .ZN(n1284) );
  aoi22d1 U1908 ( .A1(\gpio_configure[30][2] ), .A2(n1619), .B1(
        \gpio_configure[16][2] ), .B2(n1606), .ZN(n1283) );
  aoi22d1 U1909 ( .A1(\gpio_configure[8][2] ), .A2(n1578), .B1(
        \gpio_configure[13][2] ), .B2(n1582), .ZN(n1282) );
  aoi22d1 U1910 ( .A1(\gpio_configure[24][2] ), .A2(n1579), .B1(
        \gpio_configure[4][2] ), .B2(n1590), .ZN(n1289) );
  aoi22d1 U1911 ( .A1(\gpio_configure[25][2] ), .A2(n1603), .B1(
        \gpio_configure[28][2] ), .B2(n1604), .ZN(n1288) );
  aoi22d1 U1912 ( .A1(\gpio_configure[21][2] ), .A2(n1593), .B1(
        \gpio_configure[6][2] ), .B2(n1602), .ZN(n1287) );
  aoi22d1 U1913 ( .A1(\gpio_configure[26][2] ), .A2(n1592), .B1(
        \gpio_configure[5][2] ), .B2(n1618), .ZN(n1286) );
  aoi22d1 U1914 ( .A1(\gpio_configure[20][2] ), .A2(n1614), .B1(
        \gpio_configure[11][2] ), .B2(n1607), .ZN(n1293) );
  aoi22d1 U1915 ( .A1(\gpio_configure[0][2] ), .A2(n1581), .B1(
        \gpio_configure[31][2] ), .B2(n1601), .ZN(n1292) );
  aoi22d1 U1916 ( .A1(\gpio_configure[22][2] ), .A2(n1589), .B1(
        \gpio_configure[3][2] ), .B2(n1613), .ZN(n1291) );
  aoi22d1 U1917 ( .A1(\gpio_configure[19][2] ), .A2(n1577), .B1(
        \gpio_configure[2][2] ), .B2(n1583), .ZN(n1290) );
  aoi22d1 U1918 ( .A1(\gpio_configure[18][2] ), .A2(n1580), .B1(
        \gpio_configure[27][2] ), .B2(n1591), .ZN(n1297) );
  aoi22d1 U1919 ( .A1(\gpio_configure[23][2] ), .A2(n1615), .B1(
        \gpio_configure[9][2] ), .B2(n1595), .ZN(n1296) );
  aoi22d1 U1920 ( .A1(\gpio_configure[1][2] ), .A2(n1605), .B1(
        \gpio_configure[12][2] ), .B2(n1612), .ZN(n1295) );
  aoi22d1 U1921 ( .A1(\gpio_configure[10][2] ), .A2(n1616), .B1(
        \gpio_configure[14][2] ), .B2(n1594), .ZN(n1294) );
  oai22d1 U1922 ( .A1(n1303), .A2(n1630), .B1(n1302), .B2(n1628), .ZN(n1308)
         );
  inv0d0 U1923 ( .I(n1635), .ZN(n1507) );
  aoi22d1 U1924 ( .A1(\gpio_configure[33][2] ), .A2(n1633), .B1(n1632), .B2(
        serial_data_staging_2[2]), .ZN(n1305) );
  aoi22d1 U1925 ( .A1(\gpio_configure[32][2] ), .A2(n1538), .B1(
        \gpio_configure[36][2] ), .B2(n1642), .ZN(n1304) );
  oai211d1 U1926 ( .C1(n1306), .C2(n1507), .A(n1305), .B(n1304), .ZN(n1307) );
  aoi211d1 U1927 ( .C1(n1634), .C2(serial_data_staging_2[1]), .A(n1308), .B(
        n1307), .ZN(n1309) );
  oai21d1 U1928 ( .B1(n1310), .B2(n1646), .A(n1309), .ZN(n2640) );
  aoi22d1 U1929 ( .A1(\gpio_configure[26][3] ), .A2(n1592), .B1(
        \gpio_configure[8][3] ), .B2(n1578), .ZN(n1314) );
  aoi22d1 U1930 ( .A1(\gpio_configure[12][3] ), .A2(n1612), .B1(
        \gpio_configure[14][3] ), .B2(n1594), .ZN(n1313) );
  aoi22d1 U1931 ( .A1(\gpio_configure[9][3] ), .A2(n1595), .B1(
        \gpio_configure[13][3] ), .B2(n1582), .ZN(n1312) );
  aoi22d1 U1932 ( .A1(\gpio_configure[23][3] ), .A2(n1615), .B1(
        \gpio_configure[6][3] ), .B2(n1602), .ZN(n1311) );
  aoi22d1 U1933 ( .A1(\gpio_configure[29][3] ), .A2(n1617), .B1(
        \gpio_configure[16][3] ), .B2(n1606), .ZN(n1318) );
  aoi22d1 U1934 ( .A1(\gpio_configure[4][3] ), .A2(n1590), .B1(
        \gpio_configure[7][3] ), .B2(n1600), .ZN(n1317) );
  aoi22d1 U1935 ( .A1(\gpio_configure[31][3] ), .A2(n1601), .B1(
        \gpio_configure[25][3] ), .B2(n1603), .ZN(n1316) );
  aoi22d1 U1936 ( .A1(\gpio_configure[22][3] ), .A2(n1589), .B1(
        \gpio_configure[30][3] ), .B2(n1619), .ZN(n1315) );
  aoi22d1 U1937 ( .A1(\gpio_configure[18][3] ), .A2(n1580), .B1(
        \gpio_configure[19][3] ), .B2(n1577), .ZN(n1322) );
  aoi22d1 U1938 ( .A1(\gpio_configure[21][3] ), .A2(n1593), .B1(
        \gpio_configure[1][3] ), .B2(n1605), .ZN(n1321) );
  aoi22d1 U1939 ( .A1(\gpio_configure[27][3] ), .A2(n1591), .B1(
        \gpio_configure[3][3] ), .B2(n1613), .ZN(n1320) );
  aoi22d1 U1940 ( .A1(\gpio_configure[24][3] ), .A2(n1579), .B1(
        \gpio_configure[15][3] ), .B2(n1588), .ZN(n1319) );
  aoi22d1 U1941 ( .A1(\gpio_configure[0][3] ), .A2(n1581), .B1(
        \gpio_configure[28][3] ), .B2(n1604), .ZN(n1326) );
  aoi22d1 U1942 ( .A1(\gpio_configure[5][3] ), .A2(n1618), .B1(
        \gpio_configure[10][3] ), .B2(n1616), .ZN(n1325) );
  aoi22d1 U1943 ( .A1(\gpio_configure[20][3] ), .A2(n1614), .B1(
        \gpio_configure[2][3] ), .B2(n1583), .ZN(n1324) );
  aoi22d1 U1944 ( .A1(\gpio_configure[17][3] ), .A2(n1576), .B1(
        \gpio_configure[11][3] ), .B2(n1607), .ZN(n1323) );
  nr04d0 U1945 ( .A1(n1330), .A2(n1329), .A3(n1328), .A4(n1327), .ZN(n1338) );
  aoi322d1 U1946 ( .C1(n1476), .C2(serial_data_staging_2[3]), .C3(n1646), .A1(
        n1634), .A2(serial_data_staging_2[2]), .B1(n1570), .B2(
        \gpio_configure[35][3] ), .ZN(n1337) );
  oai22d1 U1947 ( .A1(n1332), .A2(n1628), .B1(n1331), .B2(n1478), .ZN(n1335)
         );
  oai22d1 U1948 ( .A1(n1333), .A2(n1638), .B1(mgmt_gpio_oeb[37]), .B2(n1507), 
        .ZN(n1334) );
  aoi211d1 U1949 ( .C1(\gpio_configure[36][3] ), .C2(n1642), .A(n1335), .B(
        n1334), .ZN(n1336) );
  oai211d1 U1950 ( .C1(n1338), .C2(n1646), .A(n1337), .B(n1336), .ZN(n2639) );
  aoi22d1 U1951 ( .A1(\gpio_configure[31][4] ), .A2(n1601), .B1(
        \gpio_configure[4][4] ), .B2(n1590), .ZN(n1342) );
  aoi22d1 U1952 ( .A1(\gpio_configure[16][4] ), .A2(n1606), .B1(
        \gpio_configure[11][4] ), .B2(n1607), .ZN(n1341) );
  aoi22d1 U1953 ( .A1(\gpio_configure[21][4] ), .A2(n1593), .B1(
        \gpio_configure[28][4] ), .B2(n1604), .ZN(n1340) );
  aoi22d1 U1954 ( .A1(\gpio_configure[0][4] ), .A2(n1581), .B1(
        \gpio_configure[13][4] ), .B2(n1582), .ZN(n1339) );
  aoi22d1 U1955 ( .A1(\gpio_configure[20][4] ), .A2(n1614), .B1(
        \gpio_configure[27][4] ), .B2(n1591), .ZN(n1346) );
  aoi22d1 U1956 ( .A1(\gpio_configure[23][4] ), .A2(n1615), .B1(
        \gpio_configure[7][4] ), .B2(n1600), .ZN(n1345) );
  aoi22d1 U1957 ( .A1(\gpio_configure[12][4] ), .A2(n1612), .B1(
        \gpio_configure[14][4] ), .B2(n1594), .ZN(n1344) );
  aoi22d1 U1958 ( .A1(\gpio_configure[17][4] ), .A2(n1576), .B1(
        \gpio_configure[10][4] ), .B2(n1616), .ZN(n1343) );
  aoi22d1 U1959 ( .A1(\gpio_configure[15][4] ), .A2(n1588), .B1(
        \gpio_configure[1][4] ), .B2(n1605), .ZN(n1350) );
  aoi22d1 U1960 ( .A1(\gpio_configure[29][4] ), .A2(n1617), .B1(
        \gpio_configure[9][4] ), .B2(n1595), .ZN(n1349) );
  aoi22d1 U1961 ( .A1(\gpio_configure[18][4] ), .A2(n1580), .B1(
        \gpio_configure[26][4] ), .B2(n1592), .ZN(n1348) );
  aoi22d1 U1962 ( .A1(\gpio_configure[24][4] ), .A2(n1579), .B1(
        \gpio_configure[5][4] ), .B2(n1618), .ZN(n1347) );
  aoi22d1 U1963 ( .A1(\gpio_configure[25][4] ), .A2(n1603), .B1(
        \gpio_configure[6][4] ), .B2(n1602), .ZN(n1354) );
  aoi22d1 U1964 ( .A1(\gpio_configure[8][4] ), .A2(n1578), .B1(
        \gpio_configure[2][4] ), .B2(n1583), .ZN(n1353) );
  aoi22d1 U1965 ( .A1(\gpio_configure[30][4] ), .A2(n1619), .B1(
        \gpio_configure[3][4] ), .B2(n1613), .ZN(n1352) );
  aoi22d1 U1966 ( .A1(\gpio_configure[22][4] ), .A2(n1589), .B1(
        \gpio_configure[19][4] ), .B2(n1577), .ZN(n1351) );
  nr04d0 U1967 ( .A1(n1358), .A2(n1357), .A3(n1356), .A4(n1355), .ZN(n1367) );
  oai22d1 U1968 ( .A1(n1360), .A2(n1507), .B1(n1359), .B2(n1478), .ZN(n1365)
         );
  aoi22d1 U1969 ( .A1(\gpio_configure[32][4] ), .A2(n1538), .B1(n1632), .B2(
        serial_data_staging_2[4]), .ZN(n1362) );
  aoi22d1 U1970 ( .A1(\gpio_configure[36][4] ), .A2(n1642), .B1(
        \gpio_configure[35][4] ), .B2(n1570), .ZN(n1361) );
  oai211d1 U1971 ( .C1(n1363), .C2(n1628), .A(n1362), .B(n1361), .ZN(n1364) );
  aoi211d1 U1972 ( .C1(n1634), .C2(serial_data_staging_2[3]), .A(n1365), .B(
        n1364), .ZN(n1366) );
  oai21d1 U1973 ( .B1(n1367), .B2(n1646), .A(n1366), .ZN(n2638) );
  aoi22d1 U1974 ( .A1(\gpio_configure[9][5] ), .A2(n1595), .B1(
        \gpio_configure[27][5] ), .B2(n1591), .ZN(n1371) );
  aoi22d1 U1975 ( .A1(\gpio_configure[10][5] ), .A2(n1616), .B1(
        \gpio_configure[15][5] ), .B2(n1588), .ZN(n1370) );
  aoi22d1 U1976 ( .A1(\gpio_configure[20][5] ), .A2(n1614), .B1(
        \gpio_configure[21][5] ), .B2(n1593), .ZN(n1369) );
  aoi22d1 U1977 ( .A1(\gpio_configure[25][5] ), .A2(n1603), .B1(
        \gpio_configure[31][5] ), .B2(n1601), .ZN(n1368) );
  aoi22d1 U1978 ( .A1(\gpio_configure[4][5] ), .A2(n1590), .B1(
        \gpio_configure[22][5] ), .B2(n1589), .ZN(n1375) );
  aoi22d1 U1979 ( .A1(\gpio_configure[14][5] ), .A2(n1594), .B1(
        \gpio_configure[18][5] ), .B2(n1580), .ZN(n1374) );
  aoi22d1 U1980 ( .A1(\gpio_configure[30][5] ), .A2(n1619), .B1(
        \gpio_configure[26][5] ), .B2(n1592), .ZN(n1373) );
  aoi22d1 U1981 ( .A1(\gpio_configure[28][5] ), .A2(n1604), .B1(
        \gpio_configure[0][5] ), .B2(n1581), .ZN(n1372) );
  aoi22d1 U1982 ( .A1(\gpio_configure[1][5] ), .A2(n1605), .B1(
        \gpio_configure[29][5] ), .B2(n1617), .ZN(n1379) );
  aoi22d1 U1983 ( .A1(\gpio_configure[5][5] ), .A2(n1618), .B1(
        \gpio_configure[7][5] ), .B2(n1600), .ZN(n1378) );
  aoi22d1 U1984 ( .A1(\gpio_configure[6][5] ), .A2(n1602), .B1(
        \gpio_configure[23][5] ), .B2(n1615), .ZN(n1377) );
  aoi22d1 U1985 ( .A1(\gpio_configure[2][5] ), .A2(n1583), .B1(
        \gpio_configure[11][5] ), .B2(n1607), .ZN(n1376) );
  aoi22d1 U1986 ( .A1(\gpio_configure[12][5] ), .A2(n1612), .B1(
        \gpio_configure[3][5] ), .B2(n1613), .ZN(n1383) );
  aoi22d1 U1987 ( .A1(\gpio_configure[8][5] ), .A2(n1578), .B1(
        \gpio_configure[19][5] ), .B2(n1577), .ZN(n1382) );
  aoi22d1 U1988 ( .A1(\gpio_configure[17][5] ), .A2(n1576), .B1(
        \gpio_configure[24][5] ), .B2(n1579), .ZN(n1381) );
  aoi22d1 U1989 ( .A1(\gpio_configure[13][5] ), .A2(n1582), .B1(
        \gpio_configure[16][5] ), .B2(n1606), .ZN(n1380) );
  nr04d0 U1990 ( .A1(n1387), .A2(n1386), .A3(n1385), .A4(n1384), .ZN(n1396) );
  aoi322d1 U1991 ( .C1(n1476), .C2(serial_data_staging_2[5]), .C3(n1646), .A1(
        \gpio_configure[36][5] ), .A2(n1642), .B1(\gpio_configure[37][5] ), 
        .B2(n1635), .ZN(n1395) );
  oai22d1 U1992 ( .A1(n1389), .A2(n1628), .B1(n1388), .B2(n1638), .ZN(n1393)
         );
  oai22d1 U1993 ( .A1(n1391), .A2(n1478), .B1(n1390), .B2(n1630), .ZN(n1392)
         );
  aoi211d1 U1994 ( .C1(n1634), .C2(serial_data_staging_2[4]), .A(n1393), .B(
        n1392), .ZN(n1394) );
  oai211d1 U1995 ( .C1(n1396), .C2(n1646), .A(n1395), .B(n1394), .ZN(n2637) );
  aoi22d1 U1996 ( .A1(\gpio_configure[8][6] ), .A2(n1578), .B1(
        \gpio_configure[28][6] ), .B2(n1604), .ZN(n1400) );
  aoi22d1 U1997 ( .A1(\gpio_configure[6][6] ), .A2(n1602), .B1(
        \gpio_configure[25][6] ), .B2(n1603), .ZN(n1399) );
  aoi22d1 U1998 ( .A1(\gpio_configure[1][6] ), .A2(n1605), .B1(
        \gpio_configure[30][6] ), .B2(n1619), .ZN(n1398) );
  aoi22d1 U1999 ( .A1(\gpio_configure[0][6] ), .A2(n1581), .B1(
        \gpio_configure[31][6] ), .B2(n1601), .ZN(n1397) );
  aoi22d1 U2000 ( .A1(\gpio_configure[21][6] ), .A2(n1593), .B1(
        \gpio_configure[17][6] ), .B2(n1576), .ZN(n1404) );
  aoi22d1 U2001 ( .A1(\gpio_configure[10][6] ), .A2(n1616), .B1(
        \gpio_configure[14][6] ), .B2(n1594), .ZN(n1403) );
  aoi22d1 U2002 ( .A1(\gpio_configure[3][6] ), .A2(n1613), .B1(
        \gpio_configure[2][6] ), .B2(n1583), .ZN(n1402) );
  aoi22d1 U2003 ( .A1(\gpio_configure[11][6] ), .A2(n1607), .B1(
        \gpio_configure[9][6] ), .B2(n1595), .ZN(n1401) );
  aoi22d1 U2004 ( .A1(\gpio_configure[12][6] ), .A2(n1612), .B1(
        \gpio_configure[29][6] ), .B2(n1617), .ZN(n1408) );
  aoi22d1 U2005 ( .A1(\gpio_configure[15][6] ), .A2(n1588), .B1(
        \gpio_configure[22][6] ), .B2(n1589), .ZN(n1407) );
  aoi22d1 U2006 ( .A1(\gpio_configure[4][6] ), .A2(n1590), .B1(
        \gpio_configure[24][6] ), .B2(n1579), .ZN(n1406) );
  aoi22d1 U2007 ( .A1(\gpio_configure[5][6] ), .A2(n1618), .B1(
        \gpio_configure[27][6] ), .B2(n1591), .ZN(n1405) );
  aoi22d1 U2008 ( .A1(\gpio_configure[13][6] ), .A2(n1582), .B1(
        \gpio_configure[7][6] ), .B2(n1600), .ZN(n1412) );
  aoi22d1 U2009 ( .A1(\gpio_configure[26][6] ), .A2(n1592), .B1(
        \gpio_configure[19][6] ), .B2(n1577), .ZN(n1411) );
  aoi22d1 U2010 ( .A1(\gpio_configure[18][6] ), .A2(n1580), .B1(
        \gpio_configure[20][6] ), .B2(n1614), .ZN(n1410) );
  aoi22d1 U2011 ( .A1(\gpio_configure[16][6] ), .A2(n1606), .B1(
        \gpio_configure[23][6] ), .B2(n1615), .ZN(n1409) );
  nr04d0 U2012 ( .A1(n1416), .A2(n1415), .A3(n1414), .A4(n1413), .ZN(n1425) );
  oai22d1 U2013 ( .A1(n1418), .A2(n1507), .B1(n1417), .B2(n1638), .ZN(n1423)
         );
  aoi22d1 U2014 ( .A1(\gpio_configure[33][6] ), .A2(n1633), .B1(n1632), .B2(
        serial_data_staging_2[6]), .ZN(n1420) );
  aoi22d1 U2015 ( .A1(\gpio_configure[35][6] ), .A2(n1570), .B1(n1634), .B2(
        serial_data_staging_2[5]), .ZN(n1419) );
  oai211d1 U2016 ( .C1(n1421), .C2(n1628), .A(n1420), .B(n1419), .ZN(n1422) );
  aoi211d1 U2017 ( .C1(\gpio_configure[36][6] ), .C2(n1642), .A(n1423), .B(
        n1422), .ZN(n1424) );
  oai21d1 U2018 ( .B1(n1425), .B2(n1646), .A(n1424), .ZN(n2636) );
  aoi22d1 U2019 ( .A1(\gpio_configure[28][7] ), .A2(n1604), .B1(
        \gpio_configure[26][7] ), .B2(n1592), .ZN(n1429) );
  aoi22d1 U2020 ( .A1(\gpio_configure[8][7] ), .A2(n1578), .B1(
        \gpio_configure[23][7] ), .B2(n1615), .ZN(n1428) );
  aoi22d1 U2021 ( .A1(\gpio_configure[14][7] ), .A2(n1594), .B1(
        \gpio_configure[17][7] ), .B2(n1576), .ZN(n1427) );
  aoi22d1 U2022 ( .A1(\gpio_configure[27][7] ), .A2(n1591), .B1(
        \gpio_configure[30][7] ), .B2(n1619), .ZN(n1426) );
  aoi22d1 U2023 ( .A1(\gpio_configure[24][7] ), .A2(n1579), .B1(
        \gpio_configure[25][7] ), .B2(n1603), .ZN(n1433) );
  aoi22d1 U2024 ( .A1(\gpio_configure[9][7] ), .A2(n1595), .B1(
        \gpio_configure[1][7] ), .B2(n1605), .ZN(n1432) );
  aoi22d1 U2025 ( .A1(\gpio_configure[5][7] ), .A2(n1618), .B1(
        \gpio_configure[19][7] ), .B2(n1577), .ZN(n1431) );
  aoi22d1 U2026 ( .A1(\gpio_configure[2][7] ), .A2(n1583), .B1(
        \gpio_configure[7][7] ), .B2(n1600), .ZN(n1430) );
  aoi22d1 U2027 ( .A1(\gpio_configure[3][7] ), .A2(n1613), .B1(
        \gpio_configure[31][7] ), .B2(n1601), .ZN(n1437) );
  aoi22d1 U2028 ( .A1(\gpio_configure[11][7] ), .A2(n1607), .B1(
        \gpio_configure[29][7] ), .B2(n1617), .ZN(n1436) );
  aoi22d1 U2029 ( .A1(\gpio_configure[10][7] ), .A2(n1616), .B1(
        \gpio_configure[20][7] ), .B2(n1614), .ZN(n1435) );
  aoi22d1 U2030 ( .A1(\gpio_configure[13][7] ), .A2(n1582), .B1(
        \gpio_configure[4][7] ), .B2(n1590), .ZN(n1434) );
  aoi22d1 U2031 ( .A1(\gpio_configure[12][7] ), .A2(n1612), .B1(
        \gpio_configure[16][7] ), .B2(n1606), .ZN(n1441) );
  aoi22d1 U2032 ( .A1(\gpio_configure[15][7] ), .A2(n1588), .B1(
        \gpio_configure[22][7] ), .B2(n1589), .ZN(n1440) );
  aoi22d1 U2033 ( .A1(\gpio_configure[21][7] ), .A2(n1593), .B1(
        \gpio_configure[0][7] ), .B2(n1581), .ZN(n1439) );
  aoi22d1 U2034 ( .A1(\gpio_configure[6][7] ), .A2(n1602), .B1(
        \gpio_configure[18][7] ), .B2(n1580), .ZN(n1438) );
  nr04d0 U2035 ( .A1(n1445), .A2(n1444), .A3(n1443), .A4(n1442), .ZN(n1455) );
  aoi322d1 U2036 ( .C1(n1672), .C2(n1446), .C3(\gpio_configure[32][7] ), .A1(
        \gpio_configure[36][7] ), .A2(n1642), .B1(serial_data_staging_2[6]), 
        .B2(n1634), .ZN(n1454) );
  oai22d1 U2037 ( .A1(n1448), .A2(n1628), .B1(n1447), .B2(n1478), .ZN(n1452)
         );
  oai22d1 U2038 ( .A1(n1450), .A2(n1507), .B1(n1449), .B2(n1630), .ZN(n1451)
         );
  aoi211d1 U2039 ( .C1(n1632), .C2(serial_data_staging_2[7]), .A(n1452), .B(
        n1451), .ZN(n1453) );
  oai211d1 U2040 ( .C1(n1455), .C2(n1646), .A(n1454), .B(n1453), .ZN(n2635) );
  aoi22d1 U2041 ( .A1(\gpio_configure[0][8] ), .A2(n1581), .B1(
        \gpio_configure[10][8] ), .B2(n1616), .ZN(n1459) );
  aoi22d1 U2042 ( .A1(\gpio_configure[3][8] ), .A2(n1613), .B1(
        \gpio_configure[16][8] ), .B2(n1606), .ZN(n1458) );
  aoi22d1 U2043 ( .A1(\gpio_configure[22][8] ), .A2(n1589), .B1(
        \gpio_configure[19][8] ), .B2(n1577), .ZN(n1457) );
  aoi22d1 U2044 ( .A1(\gpio_configure[31][8] ), .A2(n1601), .B1(
        \gpio_configure[15][8] ), .B2(n1588), .ZN(n1456) );
  aoi22d1 U2045 ( .A1(\gpio_configure[18][8] ), .A2(n1580), .B1(
        \gpio_configure[27][8] ), .B2(n1591), .ZN(n1463) );
  aoi22d1 U2046 ( .A1(\gpio_configure[20][8] ), .A2(n1614), .B1(
        \gpio_configure[11][8] ), .B2(n1607), .ZN(n1462) );
  aoi22d1 U2047 ( .A1(\gpio_configure[23][8] ), .A2(n1615), .B1(
        \gpio_configure[26][8] ), .B2(n1592), .ZN(n1461) );
  aoi22d1 U2048 ( .A1(\gpio_configure[1][8] ), .A2(n1605), .B1(
        \gpio_configure[13][8] ), .B2(n1582), .ZN(n1460) );
  aoi22d1 U2049 ( .A1(\gpio_configure[4][8] ), .A2(n1590), .B1(
        \gpio_configure[8][8] ), .B2(n1578), .ZN(n1467) );
  aoi22d1 U2050 ( .A1(\gpio_configure[24][8] ), .A2(n1579), .B1(
        \gpio_configure[14][8] ), .B2(n1594), .ZN(n1466) );
  aoi22d1 U2051 ( .A1(\gpio_configure[6][8] ), .A2(n1602), .B1(
        \gpio_configure[7][8] ), .B2(n1600), .ZN(n1465) );
  aoi22d1 U2052 ( .A1(\gpio_configure[30][8] ), .A2(n1619), .B1(
        \gpio_configure[25][8] ), .B2(n1603), .ZN(n1464) );
  aoi22d1 U2053 ( .A1(\gpio_configure[5][8] ), .A2(n1618), .B1(
        \gpio_configure[17][8] ), .B2(n1576), .ZN(n1471) );
  aoi22d1 U2054 ( .A1(\gpio_configure[29][8] ), .A2(n1617), .B1(
        \gpio_configure[9][8] ), .B2(n1595), .ZN(n1470) );
  aoi22d1 U2055 ( .A1(\gpio_configure[21][8] ), .A2(n1593), .B1(
        \gpio_configure[2][8] ), .B2(n1583), .ZN(n1469) );
  aoi22d1 U2056 ( .A1(\gpio_configure[28][8] ), .A2(n1604), .B1(
        \gpio_configure[12][8] ), .B2(n1612), .ZN(n1468) );
  aoi322d1 U2057 ( .C1(n1476), .C2(serial_data_staging_2[8]), .C3(n1646), .A1(
        n1634), .A2(serial_data_staging_2[7]), .B1(n1570), .B2(
        \gpio_configure[35][8] ), .ZN(n1485) );
  oai22d1 U2058 ( .A1(n1479), .A2(n1478), .B1(n1477), .B2(n1628), .ZN(n1483)
         );
  oai22d1 U2059 ( .A1(n1481), .A2(n1638), .B1(n1480), .B2(n1507), .ZN(n1482)
         );
  aoi211d1 U2060 ( .C1(\gpio_configure[36][8] ), .C2(n1642), .A(n1483), .B(
        n1482), .ZN(n1484) );
  oai211d1 U2061 ( .C1(n1486), .C2(n1646), .A(n1485), .B(n1484), .ZN(n2634) );
  aoi22d1 U2062 ( .A1(\gpio_configure[16][9] ), .A2(n1606), .B1(
        \gpio_configure[15][9] ), .B2(n1588), .ZN(n1490) );
  aoi22d1 U2063 ( .A1(\gpio_configure[7][9] ), .A2(n1600), .B1(
        \gpio_configure[20][9] ), .B2(n1614), .ZN(n1489) );
  aoi22d1 U2064 ( .A1(\gpio_configure[12][9] ), .A2(n1612), .B1(
        \gpio_configure[3][9] ), .B2(n1613), .ZN(n1488) );
  aoi22d1 U2065 ( .A1(\gpio_configure[6][9] ), .A2(n1602), .B1(
        \gpio_configure[18][9] ), .B2(n1580), .ZN(n1487) );
  aoi22d1 U2066 ( .A1(\gpio_configure[22][9] ), .A2(n1589), .B1(
        \gpio_configure[19][9] ), .B2(n1577), .ZN(n1494) );
  aoi22d1 U2067 ( .A1(\gpio_configure[8][9] ), .A2(n1578), .B1(
        \gpio_configure[0][9] ), .B2(n1581), .ZN(n1493) );
  aoi22d1 U2068 ( .A1(\gpio_configure[23][9] ), .A2(n1615), .B1(
        \gpio_configure[29][9] ), .B2(n1617), .ZN(n1492) );
  aoi22d1 U2069 ( .A1(\gpio_configure[2][9] ), .A2(n1583), .B1(
        \gpio_configure[1][9] ), .B2(n1605), .ZN(n1491) );
  aoi22d1 U2070 ( .A1(\gpio_configure[26][9] ), .A2(n1592), .B1(
        \gpio_configure[30][9] ), .B2(n1619), .ZN(n1498) );
  aoi22d1 U2071 ( .A1(\gpio_configure[9][9] ), .A2(n1595), .B1(
        \gpio_configure[4][9] ), .B2(n1590), .ZN(n1497) );
  aoi22d1 U2072 ( .A1(\gpio_configure[5][9] ), .A2(n1618), .B1(
        \gpio_configure[25][9] ), .B2(n1603), .ZN(n1496) );
  aoi22d1 U2073 ( .A1(\gpio_configure[13][9] ), .A2(n1582), .B1(
        \gpio_configure[28][9] ), .B2(n1604), .ZN(n1495) );
  aoi22d1 U2074 ( .A1(\gpio_configure[21][9] ), .A2(n1593), .B1(
        \gpio_configure[27][9] ), .B2(n1591), .ZN(n1502) );
  aoi22d1 U2075 ( .A1(\gpio_configure[11][9] ), .A2(n1607), .B1(
        \gpio_configure[14][9] ), .B2(n1594), .ZN(n1501) );
  aoi22d1 U2076 ( .A1(\gpio_configure[10][9] ), .A2(n1616), .B1(
        \gpio_configure[24][9] ), .B2(n1579), .ZN(n1500) );
  aoi22d1 U2077 ( .A1(\gpio_configure[17][9] ), .A2(n1576), .B1(
        \gpio_configure[31][9] ), .B2(n1601), .ZN(n1499) );
  nr04d0 U2078 ( .A1(n1506), .A2(n1505), .A3(n1504), .A4(n1503), .ZN(n1516) );
  oai22d1 U2079 ( .A1(n1509), .A2(n1630), .B1(n1508), .B2(n1507), .ZN(n1514)
         );
  aoi22d1 U2080 ( .A1(\gpio_configure[32][9] ), .A2(n1538), .B1(
        \gpio_configure[33][9] ), .B2(n1633), .ZN(n1511) );
  aoi22d1 U2081 ( .A1(\gpio_configure[36][9] ), .A2(n1642), .B1(n1634), .B2(
        serial_data_staging_2[8]), .ZN(n1510) );
  oai211d1 U2082 ( .C1(n1512), .C2(n1628), .A(n1511), .B(n1510), .ZN(n1513) );
  aoi211d1 U2083 ( .C1(n1632), .C2(serial_data_staging_2[9]), .A(n1514), .B(
        n1513), .ZN(n1515) );
  oai21d1 U2084 ( .B1(n1516), .B2(n1646), .A(n1515), .ZN(n2633) );
  aoi22d1 U2085 ( .A1(\gpio_configure[23][10] ), .A2(n1615), .B1(
        \gpio_configure[24][10] ), .B2(n1579), .ZN(n1520) );
  aoi22d1 U2086 ( .A1(\gpio_configure[15][10] ), .A2(n1588), .B1(
        \gpio_configure[11][10] ), .B2(n1607), .ZN(n1519) );
  aoi22d1 U2087 ( .A1(\gpio_configure[22][10] ), .A2(n1589), .B1(
        \gpio_configure[2][10] ), .B2(n1583), .ZN(n1518) );
  aoi22d1 U2088 ( .A1(\gpio_configure[26][10] ), .A2(n1592), .B1(
        \gpio_configure[31][10] ), .B2(n1601), .ZN(n1517) );
  aoi22d1 U2089 ( .A1(\gpio_configure[0][10] ), .A2(n1581), .B1(
        \gpio_configure[30][10] ), .B2(n1619), .ZN(n1524) );
  aoi22d1 U2090 ( .A1(\gpio_configure[29][10] ), .A2(n1617), .B1(
        \gpio_configure[14][10] ), .B2(n1594), .ZN(n1523) );
  aoi22d1 U2091 ( .A1(\gpio_configure[10][10] ), .A2(n1616), .B1(
        \gpio_configure[5][10] ), .B2(n1618), .ZN(n1522) );
  aoi22d1 U2092 ( .A1(\gpio_configure[18][10] ), .A2(n1580), .B1(
        \gpio_configure[6][10] ), .B2(n1602), .ZN(n1521) );
  aoi22d1 U2093 ( .A1(\gpio_configure[27][10] ), .A2(n1591), .B1(
        \gpio_configure[9][10] ), .B2(n1595), .ZN(n1528) );
  aoi22d1 U2094 ( .A1(\gpio_configure[13][10] ), .A2(n1582), .B1(
        \gpio_configure[17][10] ), .B2(n1576), .ZN(n1527) );
  aoi22d1 U2095 ( .A1(\gpio_configure[25][10] ), .A2(n1603), .B1(
        \gpio_configure[16][10] ), .B2(n1606), .ZN(n1526) );
  aoi22d1 U2096 ( .A1(\gpio_configure[20][10] ), .A2(n1614), .B1(
        \gpio_configure[3][10] ), .B2(n1613), .ZN(n1525) );
  aoi22d1 U2097 ( .A1(\gpio_configure[19][10] ), .A2(n1577), .B1(
        \gpio_configure[4][10] ), .B2(n1590), .ZN(n1532) );
  aoi22d1 U2098 ( .A1(\gpio_configure[1][10] ), .A2(n1605), .B1(
        \gpio_configure[28][10] ), .B2(n1604), .ZN(n1531) );
  aoi22d1 U2099 ( .A1(\gpio_configure[21][10] ), .A2(n1593), .B1(
        \gpio_configure[8][10] ), .B2(n1578), .ZN(n1530) );
  aoi22d1 U2100 ( .A1(\gpio_configure[7][10] ), .A2(n1600), .B1(
        \gpio_configure[12][10] ), .B2(n1612), .ZN(n1529) );
  nr04d0 U2101 ( .A1(n1536), .A2(n1535), .A3(n1534), .A4(n1533), .ZN(n1546) );
  aor22d1 U2102 ( .A1(\gpio_configure[37][10] ), .A2(n1635), .B1(
        \gpio_configure[34][10] ), .B2(n1537), .Z(n1544) );
  aoi22d1 U2103 ( .A1(\gpio_configure[32][10] ), .A2(n1538), .B1(
        \gpio_configure[33][10] ), .B2(n1633), .ZN(n1540) );
  aoi22d1 U2104 ( .A1(\gpio_configure[35][10] ), .A2(n1570), .B1(n1632), .B2(
        serial_data_staging_2[10]), .ZN(n1539) );
  oai211d1 U2105 ( .C1(n1542), .C2(n1541), .A(n1540), .B(n1539), .ZN(n1543) );
  aoi211d1 U2106 ( .C1(n1634), .C2(serial_data_staging_2[9]), .A(n1544), .B(
        n1543), .ZN(n1545) );
  oai21d1 U2107 ( .B1(n1546), .B2(n1646), .A(n1545), .ZN(n2632) );
  aoi22d1 U2108 ( .A1(\gpio_configure[24][11] ), .A2(n1579), .B1(
        \gpio_configure[18][11] ), .B2(n1580), .ZN(n1550) );
  aoi22d1 U2109 ( .A1(\gpio_configure[14][11] ), .A2(n1594), .B1(
        \gpio_configure[25][11] ), .B2(n1603), .ZN(n1549) );
  aoi22d1 U2110 ( .A1(\gpio_configure[8][11] ), .A2(n1578), .B1(
        \gpio_configure[28][11] ), .B2(n1604), .ZN(n1548) );
  aoi22d1 U2111 ( .A1(\gpio_configure[13][11] ), .A2(n1582), .B1(
        \gpio_configure[10][11] ), .B2(n1616), .ZN(n1547) );
  aoi22d1 U2112 ( .A1(\gpio_configure[4][11] ), .A2(n1590), .B1(
        \gpio_configure[12][11] ), .B2(n1612), .ZN(n1554) );
  aoi22d1 U2113 ( .A1(\gpio_configure[19][11] ), .A2(n1577), .B1(
        \gpio_configure[23][11] ), .B2(n1615), .ZN(n1553) );
  aoi22d1 U2114 ( .A1(\gpio_configure[16][11] ), .A2(n1606), .B1(
        \gpio_configure[7][11] ), .B2(n1600), .ZN(n1552) );
  aoi22d1 U2115 ( .A1(\gpio_configure[17][11] ), .A2(n1576), .B1(
        \gpio_configure[21][11] ), .B2(n1593), .ZN(n1551) );
  aoi22d1 U2116 ( .A1(\gpio_configure[9][11] ), .A2(n1595), .B1(
        \gpio_configure[20][11] ), .B2(n1614), .ZN(n1558) );
  aoi22d1 U2117 ( .A1(\gpio_configure[6][11] ), .A2(n1602), .B1(
        \gpio_configure[3][11] ), .B2(n1613), .ZN(n1557) );
  aoi22d1 U2118 ( .A1(\gpio_configure[1][11] ), .A2(n1605), .B1(
        \gpio_configure[27][11] ), .B2(n1591), .ZN(n1556) );
  aoi22d1 U2119 ( .A1(\gpio_configure[22][11] ), .A2(n1589), .B1(
        \gpio_configure[0][11] ), .B2(n1581), .ZN(n1555) );
  aoi22d1 U2120 ( .A1(\gpio_configure[15][11] ), .A2(n1588), .B1(
        \gpio_configure[2][11] ), .B2(n1583), .ZN(n1563) );
  aoi22d1 U2121 ( .A1(\gpio_configure[11][11] ), .A2(n1607), .B1(
        \gpio_configure[29][11] ), .B2(n1617), .ZN(n1562) );
  aoi22d1 U2122 ( .A1(\gpio_configure[5][11] ), .A2(n1618), .B1(
        \gpio_configure[31][11] ), .B2(n1601), .ZN(n1561) );
  aoi322d1 U2123 ( .C1(n1673), .C2(n1559), .C3(\gpio_configure[36][11] ), .A1(
        n1592), .A2(\gpio_configure[26][11] ), .B1(n1619), .B2(
        \gpio_configure[30][11] ), .ZN(n1560) );
  nr04d0 U2124 ( .A1(n1567), .A2(n1566), .A3(n1565), .A4(n1564), .ZN(n1575) );
  aoi22d1 U2125 ( .A1(\gpio_configure[33][11] ), .A2(n1633), .B1(n1632), .B2(
        serial_data_staging_2[11]), .ZN(n1574) );
  oai22d1 U2126 ( .A1(n1569), .A2(n1628), .B1(n1568), .B2(n1638), .ZN(n1572)
         );
  aor22d1 U2127 ( .A1(\gpio_configure[35][11] ), .A2(n1570), .B1(
        \gpio_configure[37][11] ), .B2(n1635), .Z(n1571) );
  aoi211d1 U2128 ( .C1(serial_data_staging_2[10]), .C2(n1634), .A(n1572), .B(
        n1571), .ZN(n1573) );
  oai211d1 U2129 ( .C1(n1575), .C2(n1646), .A(n1574), .B(n1573), .ZN(n2631) );
  aoi22d1 U2130 ( .A1(\gpio_configure[19][12] ), .A2(n1577), .B1(
        \gpio_configure[17][12] ), .B2(n1576), .ZN(n1587) );
  aoi22d1 U2131 ( .A1(\gpio_configure[24][12] ), .A2(n1579), .B1(
        \gpio_configure[8][12] ), .B2(n1578), .ZN(n1586) );
  aoi22d1 U2132 ( .A1(\gpio_configure[0][12] ), .A2(n1581), .B1(
        \gpio_configure[18][12] ), .B2(n1580), .ZN(n1585) );
  aoi22d1 U2133 ( .A1(\gpio_configure[2][12] ), .A2(n1583), .B1(
        \gpio_configure[13][12] ), .B2(n1582), .ZN(n1584) );
  aoi22d1 U2134 ( .A1(\gpio_configure[22][12] ), .A2(n1589), .B1(
        \gpio_configure[15][12] ), .B2(n1588), .ZN(n1599) );
  aoi22d1 U2135 ( .A1(\gpio_configure[27][12] ), .A2(n1591), .B1(
        \gpio_configure[4][12] ), .B2(n1590), .ZN(n1598) );
  aoi22d1 U2136 ( .A1(\gpio_configure[21][12] ), .A2(n1593), .B1(
        \gpio_configure[26][12] ), .B2(n1592), .ZN(n1597) );
  aoi22d1 U2137 ( .A1(\gpio_configure[9][12] ), .A2(n1595), .B1(
        \gpio_configure[14][12] ), .B2(n1594), .ZN(n1596) );
  aoi22d1 U2138 ( .A1(\gpio_configure[31][12] ), .A2(n1601), .B1(
        \gpio_configure[7][12] ), .B2(n1600), .ZN(n1611) );
  aoi22d1 U2139 ( .A1(\gpio_configure[25][12] ), .A2(n1603), .B1(
        \gpio_configure[6][12] ), .B2(n1602), .ZN(n1610) );
  aoi22d1 U2140 ( .A1(\gpio_configure[1][12] ), .A2(n1605), .B1(
        \gpio_configure[28][12] ), .B2(n1604), .ZN(n1609) );
  aoi22d1 U2141 ( .A1(\gpio_configure[11][12] ), .A2(n1607), .B1(
        \gpio_configure[16][12] ), .B2(n1606), .ZN(n1608) );
  aoi22d1 U2142 ( .A1(\gpio_configure[3][12] ), .A2(n1613), .B1(
        \gpio_configure[12][12] ), .B2(n1612), .ZN(n1623) );
  aoi22d1 U2143 ( .A1(\gpio_configure[23][12] ), .A2(n1615), .B1(
        \gpio_configure[20][12] ), .B2(n1614), .ZN(n1622) );
  aoi22d1 U2144 ( .A1(\gpio_configure[29][12] ), .A2(n1617), .B1(
        \gpio_configure[10][12] ), .B2(n1616), .ZN(n1621) );
  aoi22d1 U2145 ( .A1(\gpio_configure[30][12] ), .A2(n1619), .B1(
        \gpio_configure[5][12] ), .B2(n1618), .ZN(n1620) );
  nr04d0 U2146 ( .A1(n1627), .A2(n1626), .A3(n1625), .A4(n1624), .ZN(n1644) );
  oai22d1 U2147 ( .A1(n1631), .A2(n1630), .B1(n1629), .B2(n1628), .ZN(n1641)
         );
  aoi22d1 U2148 ( .A1(\gpio_configure[33][12] ), .A2(n1633), .B1(
        serial_data_staging_2[12]), .B2(n1632), .ZN(n1637) );
  aoi22d1 U2149 ( .A1(\gpio_configure[37][12] ), .A2(n1635), .B1(n1634), .B2(
        serial_data_staging_2[11]), .ZN(n1636) );
  oai211d1 U2150 ( .C1(n1639), .C2(n1638), .A(n1637), .B(n1636), .ZN(n1640) );
  aoi211d1 U2151 ( .C1(\gpio_configure[36][12] ), .C2(n1642), .A(n1641), .B(
        n1640), .ZN(n1643) );
  oai21d1 U2152 ( .B1(n1644), .B2(n1646), .A(n1643), .ZN(n2630) );
  oan211d1 U2153 ( .C1(n1687), .C2(serial_clock), .B(n1675), .A(n1660), .ZN(
        n1652) );
  nd02d0 U2154 ( .A1(xfer_count[1]), .A2(n1652), .ZN(n1654) );
  inv0d0 U2155 ( .I(n1654), .ZN(n1656) );
  nd02d0 U2156 ( .A1(n1646), .A2(n1645), .ZN(n1653) );
  inv0d0 U2157 ( .I(n1653), .ZN(n1647) );
  aon211d1 U2158 ( .C1(n1656), .C2(xfer_count[2]), .B(xfer_count[3]), .A(n1647), .ZN(n1648) );
  aoi31d1 U2159 ( .B1(xfer_count[3]), .B2(n1656), .B3(xfer_count[2]), .A(n1648), .ZN(n2629) );
  aoi21d1 U2160 ( .B1(n1649), .B2(xfer_state[1]), .A(xfer_count[0]), .ZN(n1650) );
  oan211d1 U2161 ( .C1(n1651), .C2(n1650), .B(n1661), .A(n1652), .ZN(n2628) );
  aoim211d1 U2162 ( .C1(xfer_count[1]), .C2(n1652), .A(n1656), .B(n1653), .ZN(
        n2627) );
  inv0d0 U2163 ( .I(xfer_count[2]), .ZN(n1655) );
  aoi221d1 U2164 ( .B1(xfer_count[2]), .B2(n1656), .C1(n1655), .C2(n1654), .A(
        n1653), .ZN(n2626) );
  inv0d0 U2165 ( .I(serial_clock_pre), .ZN(n1659) );
  nd12d0 U2166 ( .A1(xfer_count[1]), .A2(n1657), .ZN(n1665) );
  nd02d0 U2167 ( .A1(n1658), .A2(n1665), .ZN(n1663) );
  oai22d1 U2168 ( .A1(n1666), .A2(serial_clock), .B1(n1659), .B2(n1663), .ZN(
        n2625) );
  or02d0 U2169 ( .A1(n1661), .A2(n1660), .Z(n1664) );
  inv0d0 U2170 ( .I(serial_load_pre), .ZN(n1662) );
  oai22d1 U2171 ( .A1(n1665), .A2(n1664), .B1(n1663), .B2(n1662), .ZN(n2624)
         );
  nd02d0 U2172 ( .A1(n1667), .A2(n1666), .ZN(n1669) );
  oaim21d1 U2173 ( .B1(serial_busy), .B2(n1669), .A(n1668), .ZN(n2623) );
  oai21d1 U2174 ( .B1(pad_count_2[0]), .B2(n1687), .A(n1670), .ZN(n2540) );
  nd02d0 U2175 ( .A1(n1696), .A2(n1673), .ZN(n1671) );
  aon211d1 U2176 ( .C1(n1687), .C2(n1671), .B(pad_count_2[1]), .A(n1677), .ZN(
        n2539) );
  oan211d1 U2177 ( .C1(n1673), .C2(n1672), .B(xfer_state[0]), .A(xfer_state[1]), .ZN(n1674) );
  aoi22d1 U2178 ( .A1(pad_count_2[2]), .A2(n1674), .B1(n1677), .B2(n1679), 
        .ZN(n2622) );
  aon211d1 U2179 ( .C1(pad_count_2[2]), .C2(pad_count_2[3]), .B(n1675), .A(
        n1674), .ZN(n1681) );
  inv0d0 U2180 ( .I(n1681), .ZN(n1680) );
  oan211d1 U2181 ( .C1(n1679), .C2(n1677), .B(n1676), .A(n1680), .ZN(n2621) );
  or03d0 U2182 ( .A1(n1679), .A2(n1678), .A3(n1677), .Z(n1684) );
  oai21d1 U2183 ( .B1(pad_count_2[4]), .B2(n1680), .A(n1684), .ZN(n2538) );
  aoi21d1 U2184 ( .B1(xfer_state[0]), .B2(n1682), .A(n1681), .ZN(n1685) );
  aoi22d1 U2185 ( .A1(pad_count_2[5]), .A2(n1685), .B1(n1684), .B2(n1683), 
        .ZN(n2620) );
  aoi22d1 U2186 ( .A1(pad_count_1[0]), .A2(n1687), .B1(n1646), .B2(n1686), 
        .ZN(n2619) );
  aoi21d1 U2187 ( .B1(xfer_state[0]), .B2(n1688), .A(xfer_state[1]), .ZN(n1692) );
  oan211d1 U2188 ( .C1(pad_count_1[0]), .C2(n1646), .B(pad_count_1[1]), .A(
        n1692), .ZN(n2537) );
  nd02d0 U2189 ( .A1(n1696), .A2(n1690), .ZN(n1695) );
  oai21d1 U2190 ( .B1(n1692), .B2(n1691), .A(n1695), .ZN(n2618) );
  aoi21d1 U2191 ( .B1(xfer_state[0]), .B2(n1693), .A(xfer_state[1]), .ZN(n1700) );
  aoi22d1 U2192 ( .A1(pad_count_1[3]), .A2(n1700), .B1(n1695), .B2(n1694), 
        .ZN(n2617) );
  oai21d1 U2193 ( .B1(n1698), .B2(n1697), .A(n1696), .ZN(n1699) );
  oai21d1 U2194 ( .B1(pad_count_1[4]), .B2(n1700), .A(n1699), .ZN(n2536) );
  nr02d1 U2195 ( .A1(n1791), .A2(n3169), .ZN(n3239) );
  aoim22d1 U2196 ( .A1(n3239), .A2(n1702), .B1(pll_trim[12]), .B2(n3239), .Z(
        n2616) );
  nd02d0 U2197 ( .A1(n2067), .A2(n3228), .ZN(n3173) );
  inv0d0 U2198 ( .I(n3173), .ZN(n3174) );
  aoim22d1 U2199 ( .A1(n3174), .A2(n1713), .B1(pll_sel[2]), .B2(n3174), .Z(
        n2615) );
  aoim22d1 U2200 ( .A1(n3174), .A2(n1764), .B1(pll_sel[0]), .B2(n3174), .Z(
        n2614) );
  aoim22d1 U2201 ( .A1(n3174), .A2(n1712), .B1(pll90_sel[0]), .B2(n3174), .Z(
        n2612) );
  nr02d1 U2202 ( .A1(n2235), .A2(n3169), .ZN(n3129) );
  aoim22d1 U2203 ( .A1(n3129), .A2(n1702), .B1(pll_div[4]), .B2(n3129), .Z(
        n2611) );
  aoim22d1 U2204 ( .A1(n3129), .A2(n1712), .B1(pll_div[3]), .B2(n3129), .Z(
        n2610) );
  aoim22d1 U2205 ( .A1(n3129), .A2(n1714), .B1(pll_div[1]), .B2(n3129), .Z(
        n2609) );
  aoim22d1 U2206 ( .A1(n3129), .A2(n1764), .B1(pll_div[0]), .B2(n3129), .Z(
        n2608) );
  nr02d0 U2207 ( .A1(n1703), .A2(n3169), .ZN(n3180) );
  aoim22d1 U2208 ( .A1(n3180), .A2(n1764), .B1(pll_ena), .B2(n3180), .Z(n2607)
         );
  nr02d0 U2209 ( .A1(n1707), .A2(n2171), .ZN(n1706) );
  aoi211d1 U2210 ( .C1(n1706), .C2(n3181), .A(n1705), .B(n1704), .ZN(n2606) );
  nr02d0 U2211 ( .A1(n1707), .A2(n2333), .ZN(n1708) );
  mx02d1 U2212 ( .I0(reset_reg), .I1(n3268), .S(n1708), .Z(n2605) );
  nr02d0 U2213 ( .A1(n1914), .A2(n2333), .ZN(n1709) );
  aoim22d1 U2214 ( .A1(n1709), .A2(n1713), .B1(clk1_output_dest), .B2(n1709), 
        .Z(n2604) );
  aoim22d1 U2215 ( .A1(n1709), .A2(n1714), .B1(clk2_output_dest), .B2(n1709), 
        .Z(n2603) );
  aoim22d1 U2216 ( .A1(n1709), .A2(n3181), .B1(trap_output_dest), .B2(n1709), 
        .Z(n2602) );
  aoim22d1 U2217 ( .A1(n1710), .A2(n1764), .B1(irq_1_inputsrc), .B2(n1710), 
        .Z(n2601) );
  nr02d0 U2218 ( .A1(n2185), .A2(n1711), .ZN(n1715) );
  aoim22d1 U2219 ( .A1(n1715), .A2(n1764), .B1(n432), .B2(n1715), .Z(n2600) );
  aoim22d1 U2220 ( .A1(n1715), .A2(n1712), .B1(n429), .B2(n1715), .Z(n2599) );
  aoim22d1 U2221 ( .A1(n1715), .A2(n1713), .B1(n430), .B2(n1715), .Z(n2598) );
  aoim22d1 U2222 ( .A1(n1715), .A2(n1714), .B1(n431), .B2(n1715), .Z(n2597) );
  nd02d0 U2223 ( .A1(n2342), .A2(n1719), .ZN(n1758) );
  inv0d0 U2224 ( .I(mgmt_gpio_data_buf[0]), .ZN(n1720) );
  inv0d0 U2225 ( .I(n1717), .ZN(n1716) );
  aoi22d1 U2226 ( .A1(n1717), .A2(n1764), .B1(n1720), .B2(n1716), .ZN(n2596)
         );
  inv0d0 U2227 ( .I(mgmt_gpio_data_buf[1]), .ZN(n1723) );
  aoi22d1 U2228 ( .A1(n1717), .A2(n1767), .B1(n1723), .B2(n1716), .ZN(n2595)
         );
  inv0d0 U2229 ( .I(mgmt_gpio_data_buf[2]), .ZN(n1725) );
  aoi22d1 U2230 ( .A1(n1717), .A2(n873), .B1(n1725), .B2(n1716), .ZN(n2594) );
  inv0d0 U2231 ( .I(mgmt_gpio_data_buf[3]), .ZN(n1727) );
  aoi22d1 U2232 ( .A1(n1717), .A2(n1772), .B1(n1727), .B2(n1716), .ZN(n2593)
         );
  inv0d0 U2233 ( .I(mgmt_gpio_data_buf[4]), .ZN(n1729) );
  aoi22d1 U2234 ( .A1(n1717), .A2(n1775), .B1(n1729), .B2(n1716), .ZN(n2592)
         );
  inv0d0 U2235 ( .I(mgmt_gpio_data_buf[5]), .ZN(n1731) );
  aoi22d1 U2236 ( .A1(n1717), .A2(n1779), .B1(n1731), .B2(n1716), .ZN(n2591)
         );
  inv0d0 U2237 ( .I(mgmt_gpio_data_buf[6]), .ZN(n1733) );
  aoi22d1 U2238 ( .A1(n1717), .A2(n1782), .B1(n1733), .B2(n1716), .ZN(n2590)
         );
  inv0d0 U2239 ( .I(mgmt_gpio_data_buf[7]), .ZN(n1737) );
  aoi22d1 U2240 ( .A1(n1717), .A2(n1786), .B1(n1737), .B2(n1716), .ZN(n2589)
         );
  nd02d0 U2241 ( .A1(n1719), .A2(n1718), .ZN(n1762) );
  inv0d0 U2242 ( .I(n2211), .ZN(n2247) );
  nr02d0 U2243 ( .A1(n1790), .A2(n2247), .ZN(n2285) );
  nd12d0 U2244 ( .A1(n1758), .A2(n2285), .ZN(n1785) );
  oai21d1 U2245 ( .B1(n633), .B2(n1762), .A(n1778), .ZN(n1735) );
  nd02d0 U2246 ( .A1(n2284), .A2(n1735), .ZN(n1736) );
  oai222d1 U2247 ( .A1(n1721), .A2(n1735), .B1(n1736), .B2(n1764), .C1(n1720), 
        .C2(n1785), .ZN(n2588) );
  oai222d1 U2248 ( .A1(n1723), .A2(n1778), .B1(n1736), .B2(n1767), .C1(n1735), 
        .C2(n1722), .ZN(n2587) );
  inv0d0 U2249 ( .I(mgmt_gpio_out[2]), .ZN(n1724) );
  oai222d1 U2250 ( .A1(n1725), .A2(n1778), .B1(n1736), .B2(n849), .C1(n1735), 
        .C2(n1724), .ZN(n2586) );
  inv0d0 U2251 ( .I(mgmt_gpio_out[3]), .ZN(n1726) );
  oai222d1 U2252 ( .A1(n1727), .A2(n1778), .B1(n1736), .B2(n1772), .C1(n1735), 
        .C2(n1726), .ZN(n2585) );
  inv0d0 U2253 ( .I(mgmt_gpio_out[4]), .ZN(n1728) );
  oai222d1 U2254 ( .A1(n1729), .A2(n1778), .B1(n1736), .B2(n1775), .C1(n1735), 
        .C2(n1728), .ZN(n2584) );
  inv0d0 U2255 ( .I(mgmt_gpio_out[5]), .ZN(n1730) );
  oai222d1 U2256 ( .A1(n1731), .A2(n1778), .B1(n1736), .B2(n1779), .C1(n1735), 
        .C2(n1730), .ZN(n2583) );
  inv0d0 U2257 ( .I(mgmt_gpio_data_6), .ZN(n1732) );
  oai222d1 U2258 ( .A1(n1733), .A2(n1778), .B1(n1736), .B2(n1782), .C1(n1735), 
        .C2(n1732), .ZN(n2582) );
  inv0d0 U2259 ( .I(mgmt_gpio_out[7]), .ZN(n1734) );
  oai222d1 U2260 ( .A1(n1737), .A2(n1778), .B1(n1736), .B2(n1786), .C1(n1735), 
        .C2(n1734), .ZN(n2581) );
  inv0d0 U2261 ( .I(mgmt_gpio_data_buf[8]), .ZN(n1741) );
  inv0d0 U2262 ( .I(n1739), .ZN(n1738) );
  aoi22d1 U2263 ( .A1(n1739), .A2(n1764), .B1(n1741), .B2(n1738), .ZN(n2580)
         );
  inv0d0 U2264 ( .I(mgmt_gpio_data_buf[9]), .ZN(n1743) );
  aoi22d1 U2265 ( .A1(n1739), .A2(n1767), .B1(n1743), .B2(n1738), .ZN(n2579)
         );
  inv0d0 U2266 ( .I(mgmt_gpio_data_buf[10]), .ZN(n1745) );
  aoi22d1 U2267 ( .A1(n1739), .A2(n849), .B1(n1745), .B2(n1738), .ZN(n2578) );
  inv0d0 U2268 ( .I(mgmt_gpio_data_buf[11]), .ZN(n1746) );
  aoi22d1 U2269 ( .A1(n1739), .A2(n1772), .B1(n1746), .B2(n1738), .ZN(n2577)
         );
  inv0d0 U2270 ( .I(mgmt_gpio_data_buf[12]), .ZN(n1748) );
  aoi22d1 U2271 ( .A1(n1739), .A2(n1775), .B1(n1748), .B2(n1738), .ZN(n2576)
         );
  inv0d0 U2272 ( .I(mgmt_gpio_data_buf[13]), .ZN(n1750) );
  aoi22d1 U2273 ( .A1(n1739), .A2(n1779), .B1(n1750), .B2(n1738), .ZN(n2575)
         );
  inv0d0 U2274 ( .I(mgmt_gpio_data_buf[14]), .ZN(n1753) );
  aoi22d1 U2275 ( .A1(n1739), .A2(n1782), .B1(n1753), .B2(n1738), .ZN(n2574)
         );
  inv0d0 U2276 ( .I(mgmt_gpio_data_buf[15]), .ZN(n1757) );
  aoi22d1 U2277 ( .A1(n1739), .A2(n1786), .B1(n1757), .B2(n1738), .ZN(n2573)
         );
  oai21d1 U2278 ( .B1(n1740), .B2(n1762), .A(n1778), .ZN(n1754) );
  nd02d0 U2279 ( .A1(n620), .A2(n1754), .ZN(n1756) );
  oai222d1 U2280 ( .A1(n1742), .A2(n1754), .B1(n1756), .B2(n1764), .C1(n1785), 
        .C2(n1741), .ZN(n2572) );
  oai222d1 U2281 ( .A1(n2319), .A2(n1754), .B1(n1756), .B2(n1767), .C1(n1743), 
        .C2(n1778), .ZN(n2571) );
  oai222d1 U2282 ( .A1(n1745), .A2(n1778), .B1(n1756), .B2(n849), .C1(n1744), 
        .C2(n1754), .ZN(n2570) );
  inv0d0 U2283 ( .I(mgmt_gpio_out[11]), .ZN(n1747) );
  oai222d1 U2284 ( .A1(n1747), .A2(n1754), .B1(n1756), .B2(n1772), .C1(n1746), 
        .C2(n1778), .ZN(n2569) );
  inv0d0 U2285 ( .I(mgmt_gpio_out[12]), .ZN(n1749) );
  oai222d1 U2286 ( .A1(n1749), .A2(n1754), .B1(n1756), .B2(n1775), .C1(n1748), 
        .C2(n1778), .ZN(n2568) );
  oai222d1 U2287 ( .A1(n1751), .A2(n1754), .B1(n1756), .B2(n1779), .C1(n1750), 
        .C2(n1778), .ZN(n2567) );
  inv0d0 U2288 ( .I(mgmt_gpio_data_14), .ZN(n1752) );
  oai222d1 U2289 ( .A1(n1753), .A2(n1778), .B1(n1756), .B2(n1782), .C1(n1752), 
        .C2(n1754), .ZN(n2566) );
  inv0d0 U2290 ( .I(mgmt_gpio_data_15), .ZN(n1755) );
  oai222d1 U2291 ( .A1(n1757), .A2(n1778), .B1(n1756), .B2(n1786), .C1(n1755), 
        .C2(n1754), .ZN(n2565) );
  nr02d0 U2292 ( .A1(n1790), .A2(n2054), .ZN(n2283) );
  nd12d0 U2293 ( .A1(n1758), .A2(n2283), .ZN(n1760) );
  inv0d0 U2294 ( .I(n1760), .ZN(n1761) );
  inv0d0 U2295 ( .I(mgmt_gpio_data_buf[16]), .ZN(n1765) );
  aoi22d1 U2296 ( .A1(n1761), .A2(n1764), .B1(n1765), .B2(n1760), .ZN(n2564)
         );
  inv0d0 U2297 ( .I(mgmt_gpio_data_buf[17]), .ZN(n1766) );
  aoi22d1 U2298 ( .A1(n1761), .A2(n1759), .B1(n1766), .B2(n1760), .ZN(n2563)
         );
  inv0d0 U2299 ( .I(mgmt_gpio_data_buf[18]), .ZN(n1769) );
  aoi22d1 U2300 ( .A1(n1761), .A2(n849), .B1(n1769), .B2(n1760), .ZN(n2562) );
  inv0d0 U2301 ( .I(mgmt_gpio_data_buf[19]), .ZN(n1771) );
  aoi22d1 U2302 ( .A1(n1761), .A2(n1772), .B1(n1771), .B2(n1760), .ZN(n2561)
         );
  inv0d0 U2303 ( .I(mgmt_gpio_data_buf[20]), .ZN(n1774) );
  aoi22d1 U2304 ( .A1(n1761), .A2(n1775), .B1(n1774), .B2(n1760), .ZN(n2560)
         );
  inv0d0 U2305 ( .I(mgmt_gpio_data_buf[21]), .ZN(n1777) );
  aoi22d1 U2306 ( .A1(n1761), .A2(n1779), .B1(n1777), .B2(n1760), .ZN(n2559)
         );
  inv0d0 U2307 ( .I(mgmt_gpio_data_buf[22]), .ZN(n1781) );
  aoi22d1 U2308 ( .A1(n1761), .A2(n1782), .B1(n1781), .B2(n1760), .ZN(n2558)
         );
  inv0d0 U2309 ( .I(mgmt_gpio_data_buf[23]), .ZN(n1784) );
  aoi22d1 U2310 ( .A1(n1761), .A2(n1786), .B1(n1784), .B2(n1760), .ZN(n2557)
         );
  nd12d0 U2311 ( .A1(n1762), .A2(n2283), .ZN(n1787) );
  inv0d0 U2312 ( .I(mgmt_gpio_out[16]), .ZN(n1763) );
  nd02d0 U2313 ( .A1(n1778), .A2(n1787), .ZN(n1789) );
  oai222d1 U2314 ( .A1(n1765), .A2(n1778), .B1(n1787), .B2(n1764), .C1(n1763), 
        .C2(n1789), .ZN(n2556) );
  inv0d0 U2315 ( .I(mgmt_gpio_out[17]), .ZN(n1768) );
  oai222d1 U2316 ( .A1(n1789), .A2(n1768), .B1(n1787), .B2(n1767), .C1(n1785), 
        .C2(n1766), .ZN(n2555) );
  inv0d0 U2317 ( .I(mgmt_gpio_out[18]), .ZN(n1770) );
  oai222d1 U2318 ( .A1(n1789), .A2(n1770), .B1(n1787), .B2(n873), .C1(n1785), 
        .C2(n1769), .ZN(n2554) );
  inv0d0 U2319 ( .I(mgmt_gpio_out[19]), .ZN(n1773) );
  oai222d1 U2320 ( .A1(n1789), .A2(n1773), .B1(n1787), .B2(n1772), .C1(n1785), 
        .C2(n1771), .ZN(n2553) );
  inv0d0 U2321 ( .I(mgmt_gpio_out[20]), .ZN(n1776) );
  oai222d1 U2322 ( .A1(n1789), .A2(n1776), .B1(n1787), .B2(n1775), .C1(n1785), 
        .C2(n1774), .ZN(n2552) );
  inv0d0 U2323 ( .I(mgmt_gpio_out[21]), .ZN(n1780) );
  oai222d1 U2324 ( .A1(n1789), .A2(n1780), .B1(n1787), .B2(n1779), .C1(n1778), 
        .C2(n1777), .ZN(n2551) );
  inv0d0 U2325 ( .I(mgmt_gpio_out[22]), .ZN(n1783) );
  oai222d1 U2326 ( .A1(n1789), .A2(n1783), .B1(n1787), .B2(n1782), .C1(n1785), 
        .C2(n1781), .ZN(n2550) );
  inv0d0 U2327 ( .I(mgmt_gpio_out[23]), .ZN(n1788) );
  oai222d1 U2328 ( .A1(n1789), .A2(n1788), .B1(n1787), .B2(n1786), .C1(n1785), 
        .C2(n1784), .ZN(n2549) );
  inv0d0 U2329 ( .I(\hkspi/ldata[0] ), .ZN(n1933) );
  aoi22d1 U2330 ( .A1(n2276), .A2(\gpio_configure[31][0] ), .B1(n2258), .B2(
        \gpio_configure[30][0] ), .ZN(n1806) );
  aoi22d1 U2331 ( .A1(n2252), .A2(\gpio_configure[20][0] ), .B1(n2241), .B2(
        irq[0]), .ZN(n1805) );
  inv0d1 U2332 ( .I(n1790), .ZN(n2269) );
  aoi22d1 U2333 ( .A1(n2269), .A2(\gpio_configure[22][0] ), .B1(n2225), .B2(
        \gpio_configure[19][0] ), .ZN(n1794) );
  aoi22d1 U2334 ( .A1(n2266), .A2(\gpio_configure[29][0] ), .B1(n2263), .B2(
        \gpio_configure[26][0] ), .ZN(n1793) );
  inv0d1 U2335 ( .I(n1791), .ZN(n3229) );
  aoi22d1 U2336 ( .A1(n3229), .A2(pll_trim[8]), .B1(n2265), .B2(
        \gpio_configure[28][0] ), .ZN(n1792) );
  aoi211d1 U2337 ( .C1(n2001), .C2(\gpio_configure[21][0] ), .A(n844), .B(
        n1795), .ZN(n1804) );
  aoi22d1 U2338 ( .A1(n2253), .A2(\gpio_configure[27][0] ), .B1(n2067), .B2(
        pll_trim[24]), .ZN(n1796) );
  oaim21d1 U2339 ( .B1(n2195), .B2(\gpio_configure[23][0] ), .A(n1796), .ZN(
        n1802) );
  inv0d1 U2340 ( .I(n2235), .ZN(n2206) );
  aoi22d1 U2341 ( .A1(n2206), .A2(pll_div[0]), .B1(n2255), .B2(
        \gpio_configure[25][0] ), .ZN(n1800) );
  aoi22d1 U2342 ( .A1(n2256), .A2(\gpio_configure[0][0] ), .B1(n2041), .B2(
        \gpio_configure[18][0] ), .ZN(n1799) );
  aoi22d1 U2343 ( .A1(n2223), .A2(irq_1_inputsrc), .B1(n2264), .B2(
        \gpio_configure[24][0] ), .ZN(n1798) );
  aoi211d1 U2344 ( .C1(n2254), .C2(\gpio_configure[32][0] ), .A(n1802), .B(
        n1801), .ZN(n1803) );
  buffd1 U2345 ( .I(n2067), .Z(n2237) );
  aoi22d1 U2346 ( .A1(n2264), .A2(\gpio_configure[25][8] ), .B1(n2237), .B2(
        pll_sel[0]), .ZN(n1810) );
  aoi22d1 U2347 ( .A1(n2253), .A2(\gpio_configure[28][8] ), .B1(n2041), .B2(
        \gpio_configure[19][8] ), .ZN(n1809) );
  aoi22d1 U2348 ( .A1(n2269), .A2(\gpio_configure[23][8] ), .B1(n2258), .B2(
        \gpio_configure[31][8] ), .ZN(n1808) );
  aoi22d1 U2349 ( .A1(n2281), .A2(pll_trim[0]), .B1(n2225), .B2(
        \gpio_configure[20][8] ), .ZN(n1807) );
  aoi22d1 U2350 ( .A1(n2252), .A2(\gpio_configure[21][8] ), .B1(n2268), .B2(
        \gpio_configure[24][8] ), .ZN(n1814) );
  aoi22d1 U2351 ( .A1(n2265), .A2(\gpio_configure[29][8] ), .B1(n2255), .B2(
        \gpio_configure[26][8] ), .ZN(n1813) );
  aoi22d1 U2352 ( .A1(n2256), .A2(\gpio_configure[1][8] ), .B1(n858), .B2(
        pll_bypass), .ZN(n1812) );
  aoi22d1 U2353 ( .A1(n2276), .A2(\gpio_configure[32][8] ), .B1(n2223), .B2(
        \gpio_configure[0][8] ), .ZN(n1811) );
  aoi22d1 U2354 ( .A1(n844), .A2(trap_output_dest), .B1(n2241), .B2(reset), 
        .ZN(n1820) );
  inv0d1 U2355 ( .I(n1815), .ZN(n2231) );
  aoi22d1 U2356 ( .A1(n2231), .A2(\gpio_configure[18][8] ), .B1(n2254), .B2(
        \gpio_configure[33][8] ), .ZN(n1819) );
  aoi22d1 U2357 ( .A1(n2142), .A2(serial_busy), .B1(n2266), .B2(
        \gpio_configure[30][8] ), .ZN(n1818) );
  aor22d1 U2358 ( .A1(n3229), .A2(pll_trim[16]), .B1(n2001), .B2(
        \gpio_configure[22][8] ), .Z(n1816) );
  aoi211d1 U2359 ( .C1(n2263), .C2(\gpio_configure[27][8] ), .A(n2238), .B(
        n1816), .ZN(n1817) );
  nr03d0 U2360 ( .A1(n1823), .A2(n1822), .A3(n1821), .ZN(n1856) );
  aoi22d1 U2361 ( .A1(n858), .A2(\gpio_configure[6][8] ), .B1(n2238), .B2(
        \gpio_configure[3][8] ), .ZN(n1827) );
  aoi22d1 U2362 ( .A1(n2256), .A2(\gpio_configure[17][8] ), .B1(n2241), .B2(
        \gpio_configure[7][8] ), .ZN(n1826) );
  aoi22d1 U2363 ( .A1(n2068), .A2(\gpio_configure[16][8] ), .B1(n2041), .B2(
        \gpio_configure[35][8] ), .ZN(n1825) );
  aoi22d1 U2364 ( .A1(n2267), .A2(\gpio_configure[34][8] ), .B1(n2094), .B2(
        \gpio_configure[36][8] ), .ZN(n1824) );
  aoi22d1 U2365 ( .A1(n2252), .A2(\gpio_configure[37][8] ), .B1(n2142), .B2(
        \gpio_configure[11][8] ), .ZN(n1831) );
  aoi22d1 U2366 ( .A1(n3229), .A2(\gpio_configure[9][8] ), .B1(n2240), .B2(
        \gpio_configure[13][8] ), .ZN(n1830) );
  aoi22d1 U2367 ( .A1(n2237), .A2(\gpio_configure[10][8] ), .B1(n2236), .B2(
        \gpio_configure[14][8] ), .ZN(n1829) );
  aoi22d1 U2368 ( .A1(n2242), .A2(\gpio_configure[2][8] ), .B1(n2001), .B2(
        mgmt_gpio_in[32]), .ZN(n1828) );
  aoi22d1 U2369 ( .A1(n2269), .A2(mgmt_gpio_in[16]), .B1(n2222), .B2(
        \gpio_configure[5][8] ), .ZN(n1835) );
  aoi22d1 U2370 ( .A1(n2230), .A2(\gpio_configure[4][8] ), .B1(n2224), .B2(
        \gpio_configure[12][8] ), .ZN(n1834) );
  aoi22d1 U2371 ( .A1(n2205), .A2(\gpio_configure[8][8] ), .B1(n2268), .B2(
        mgmt_gpio_in[0]), .ZN(n1833) );
  aoi22d1 U2372 ( .A1(n844), .A2(\gpio_configure[15][8] ), .B1(n2264), .B2(
        hkspi_disable), .ZN(n1832) );
  oai31d1 U2373 ( .B1(n1838), .B2(n1837), .B3(n1836), .A(n2131), .ZN(n1855) );
  aoi22d1 U2374 ( .A1(n2195), .A2(mgmt_gpio_in[8]), .B1(n2238), .B2(
        \gpio_configure[2][0] ), .ZN(n1842) );
  aoi22d1 U2375 ( .A1(n2242), .A2(\gpio_configure[1][0] ), .B1(n2067), .B2(
        \gpio_configure[9][0] ), .ZN(n1841) );
  aoi22d1 U2376 ( .A1(n2256), .A2(\gpio_configure[16][0] ), .B1(n2222), .B2(
        \gpio_configure[4][0] ), .ZN(n1840) );
  aoi22d1 U2377 ( .A1(n2267), .A2(\gpio_configure[33][0] ), .B1(n2269), .B2(
        mgmt_gpio_in[24]), .ZN(n1839) );
  aoi22d1 U2378 ( .A1(n844), .A2(\gpio_configure[14][0] ), .B1(n2225), .B2(
        \gpio_configure[35][0] ), .ZN(n1846) );
  aoi22d1 U2379 ( .A1(n2252), .A2(\gpio_configure[36][0] ), .B1(n2041), .B2(
        \gpio_configure[34][0] ), .ZN(n1845) );
  aoi22d1 U2380 ( .A1(n2205), .A2(\gpio_configure[7][0] ), .B1(n858), .B2(
        \gpio_configure[5][0] ), .ZN(n1844) );
  aoi22d1 U2381 ( .A1(n3229), .A2(\gpio_configure[8][0] ), .B1(n2236), .B2(
        \gpio_configure[13][0] ), .ZN(n1843) );
  aoi22d1 U2382 ( .A1(n2001), .A2(\gpio_configure[37][0] ), .B1(n2241), .B2(
        \gpio_configure[6][0] ), .ZN(n1850) );
  aoi22d1 U2383 ( .A1(n2068), .A2(\gpio_configure[15][0] ), .B1(n2230), .B2(
        \gpio_configure[3][0] ), .ZN(n1849) );
  aoi22d1 U2384 ( .A1(n2142), .A2(\gpio_configure[10][0] ), .B1(n2224), .B2(
        \gpio_configure[11][0] ), .ZN(n1848) );
  aoi22d1 U2385 ( .A1(n2264), .A2(n432), .B1(n2240), .B2(
        \gpio_configure[12][0] ), .ZN(n1847) );
  oai31d1 U2386 ( .B1(n1853), .B2(n1852), .B3(n1851), .A(n2211), .ZN(n1854) );
  oai211d1 U2387 ( .C1(n1856), .C2(n2288), .A(n1855), .B(n1854), .ZN(n1857) );
  aon211d1 U2388 ( .C1(n2220), .C2(n1858), .B(n1857), .A(n2290), .ZN(n3283) );
  nr03d0 U2389 ( .A1(\hkspi/count[2] ), .A2(\hkspi/count[1] ), .A3(
        \hkspi/count[0] ), .ZN(n2305) );
  nd02d0 U2390 ( .A1(n2305), .A2(n2296), .ZN(n2298) );
  oai22d1 U2391 ( .A1(n2296), .A2(n1933), .B1(n3283), .B2(n2298), .ZN(n2548)
         );
  aoi22d1 U2392 ( .A1(n844), .A2(\gpio_configure[14][1] ), .B1(n2200), .B2(
        mgmt_gpio_in[25]), .ZN(n1862) );
  aoi22d1 U2393 ( .A1(n3229), .A2(\gpio_configure[8][1] ), .B1(n2267), .B2(
        \gpio_configure[33][1] ), .ZN(n1861) );
  aoi22d1 U2394 ( .A1(n2268), .A2(mgmt_gpio_in[9]), .B1(n2241), .B2(
        \gpio_configure[6][1] ), .ZN(n1860) );
  aoi22d1 U2395 ( .A1(n2252), .A2(\gpio_configure[36][1] ), .B1(n2281), .B2(
        \gpio_configure[7][1] ), .ZN(n1859) );
  inv0d1 U2396 ( .I(n1863), .ZN(n2251) );
  inv0d1 U2397 ( .I(n2072), .ZN(n2257) );
  aoi22d1 U2398 ( .A1(n2251), .A2(\gpio_configure[37][1] ), .B1(n2257), .B2(
        \gpio_configure[34][1] ), .ZN(n1867) );
  aoi22d1 U2399 ( .A1(n2242), .A2(\gpio_configure[1][1] ), .B1(n2236), .B2(
        \gpio_configure[13][1] ), .ZN(n1866) );
  aoi22d1 U2400 ( .A1(n2264), .A2(n431), .B1(n2222), .B2(
        \gpio_configure[4][1] ), .ZN(n1865) );
  aoi22d1 U2401 ( .A1(n2237), .A2(\gpio_configure[9][1] ), .B1(n2238), .B2(
        \gpio_configure[2][1] ), .ZN(n1864) );
  aoi22d1 U2402 ( .A1(n858), .A2(\gpio_configure[5][1] ), .B1(n2230), .B2(
        \gpio_configure[3][1] ), .ZN(n1871) );
  aoi22d1 U2403 ( .A1(n2256), .A2(\gpio_configure[16][1] ), .B1(n2223), .B2(
        \gpio_configure[15][1] ), .ZN(n1870) );
  aoi22d1 U2404 ( .A1(n2206), .A2(\gpio_configure[10][1] ), .B1(n2224), .B2(
        \gpio_configure[11][1] ), .ZN(n1869) );
  aoi22d1 U2405 ( .A1(n2225), .A2(\gpio_configure[35][1] ), .B1(n2240), .B2(
        \gpio_configure[12][1] ), .ZN(n1868) );
  nr03d0 U2406 ( .A1(n1874), .A2(n1873), .A3(n1872), .ZN(n1894) );
  oai22d1 U2407 ( .A1(n1877), .A2(n1876), .B1(n2072), .B2(n1875), .ZN(n1892)
         );
  aoi22d1 U2408 ( .A1(n844), .A2(clk2_output_dest), .B1(n2266), .B2(
        \gpio_configure[30][9] ), .ZN(n1879) );
  aoi22d1 U2409 ( .A1(n2276), .A2(\gpio_configure[32][9] ), .B1(n2264), .B2(
        \gpio_configure[25][9] ), .ZN(n1878) );
  oai211d1 U2410 ( .C1(n2164), .C2(n1880), .A(n1879), .B(n1878), .ZN(n1891) );
  aoi22d1 U2411 ( .A1(n2252), .A2(\gpio_configure[21][9] ), .B1(n2237), .B2(
        pll_sel[1]), .ZN(n1884) );
  aoi22d1 U2412 ( .A1(n2265), .A2(\gpio_configure[29][9] ), .B1(n2094), .B2(
        \gpio_configure[20][9] ), .ZN(n1883) );
  aoi22d1 U2413 ( .A1(n2253), .A2(\gpio_configure[28][9] ), .B1(n2263), .B2(
        \gpio_configure[27][9] ), .ZN(n1882) );
  aoi22d1 U2414 ( .A1(n2254), .A2(\gpio_configure[33][9] ), .B1(n2258), .B2(
        \gpio_configure[31][9] ), .ZN(n1881) );
  aoi22d1 U2415 ( .A1(n2255), .A2(\gpio_configure[26][9] ), .B1(n2281), .B2(
        pll_trim[1]), .ZN(n1888) );
  aoi22d1 U2416 ( .A1(n2206), .A2(serial_bb_enable), .B1(n2001), .B2(
        \gpio_configure[22][9] ), .ZN(n1887) );
  aoi22d1 U2417 ( .A1(n3229), .A2(pll_trim[17]), .B1(n2200), .B2(
        \gpio_configure[23][9] ), .ZN(n1886) );
  aoi22d1 U2418 ( .A1(n2231), .A2(\gpio_configure[18][9] ), .B1(n2195), .B2(
        \gpio_configure[24][9] ), .ZN(n1885) );
  nr04d0 U2419 ( .A1(n1892), .A2(n1891), .A3(n1890), .A4(n1889), .ZN(n1893) );
  oai22d1 U2420 ( .A1(n1894), .A2(n2247), .B1(n1893), .B2(n2288), .ZN(n1932)
         );
  oai22d1 U2421 ( .A1(n1898), .A2(n1897), .B1(n1896), .B2(n1895), .ZN(n1913)
         );
  aoi22d1 U2422 ( .A1(n2256), .A2(\gpio_configure[17][9] ), .B1(n2225), .B2(
        \gpio_configure[36][9] ), .ZN(n1900) );
  aoi22d1 U2423 ( .A1(n2206), .A2(\gpio_configure[11][9] ), .B1(n2001), .B2(
        mgmt_gpio_in[33]), .ZN(n1899) );
  oai211d1 U2424 ( .C1(n2334), .C2(n1901), .A(n1900), .B(n1899), .ZN(n1912) );
  aoi22d1 U2425 ( .A1(n2231), .A2(\gpio_configure[34][9] ), .B1(n2257), .B2(
        \gpio_configure[35][9] ), .ZN(n1905) );
  aoi22d1 U2426 ( .A1(n844), .A2(\gpio_configure[15][9] ), .B1(n2268), .B2(
        mgmt_gpio_in[1]), .ZN(n1904) );
  aoi22d1 U2427 ( .A1(n2240), .A2(\gpio_configure[13][9] ), .B1(n2230), .B2(
        \gpio_configure[4][9] ), .ZN(n1903) );
  aoi22d1 U2428 ( .A1(n2252), .A2(\gpio_configure[37][9] ), .B1(n2241), .B2(
        \gpio_configure[7][9] ), .ZN(n1902) );
  aoi22d1 U2429 ( .A1(n2237), .A2(\gpio_configure[10][9] ), .B1(n858), .B2(
        \gpio_configure[6][9] ), .ZN(n1909) );
  aoi22d1 U2430 ( .A1(n2223), .A2(\gpio_configure[16][9] ), .B1(n2269), .B2(
        mgmt_gpio_in[17]), .ZN(n1908) );
  aoi22d1 U2431 ( .A1(n2242), .A2(\gpio_configure[2][9] ), .B1(n2238), .B2(
        \gpio_configure[3][9] ), .ZN(n1907) );
  aoi22d1 U2432 ( .A1(n2282), .A2(\gpio_configure[9][9] ), .B1(n2224), .B2(
        \gpio_configure[12][9] ), .ZN(n1906) );
  nr04d0 U2433 ( .A1(n1913), .A2(n1912), .A3(n1911), .A4(n1910), .ZN(n1930) );
  nd02d0 U2434 ( .A1(n1914), .A2(n2150), .ZN(n1953) );
  aoi22d1 U2435 ( .A1(n2256), .A2(\gpio_configure[0][1] ), .B1(n2237), .B2(
        pll_trim[25]), .ZN(n1917) );
  aoi22d1 U2436 ( .A1(n2252), .A2(\gpio_configure[20][1] ), .B1(n2001), .B2(
        \gpio_configure[21][1] ), .ZN(n1916) );
  aoi22d1 U2437 ( .A1(n2231), .A2(\gpio_configure[17][1] ), .B1(n2255), .B2(
        \gpio_configure[25][1] ), .ZN(n1915) );
  aoi22d1 U2438 ( .A1(n2265), .A2(\gpio_configure[28][1] ), .B1(n2195), .B2(
        \gpio_configure[23][1] ), .ZN(n1921) );
  aoi22d1 U2439 ( .A1(n2269), .A2(\gpio_configure[22][1] ), .B1(n2253), .B2(
        \gpio_configure[27][1] ), .ZN(n1920) );
  aoi22d1 U2440 ( .A1(n2276), .A2(\gpio_configure[31][1] ), .B1(n2263), .B2(
        \gpio_configure[26][1] ), .ZN(n1919) );
  aoi22d1 U2441 ( .A1(n3229), .A2(pll_trim[9]), .B1(n2266), .B2(
        \gpio_configure[29][1] ), .ZN(n1918) );
  aoi22d1 U2442 ( .A1(n2264), .A2(\gpio_configure[24][1] ), .B1(n2258), .B2(
        \gpio_configure[30][1] ), .ZN(n1925) );
  aoi22d1 U2443 ( .A1(n2225), .A2(\gpio_configure[19][1] ), .B1(n2041), .B2(
        \gpio_configure[18][1] ), .ZN(n1924) );
  aoi22d1 U2444 ( .A1(n2206), .A2(pll_div[1]), .B1(n2223), .B2(irq_2_inputsrc), 
        .ZN(n1923) );
  aoi22d1 U2445 ( .A1(n2254), .A2(\gpio_configure[32][1] ), .B1(n858), .B2(
        pll_dco_ena), .ZN(n1922) );
  oai22d1 U2446 ( .A1(n1930), .A2(n2054), .B1(n1929), .B2(n2277), .ZN(n1931)
         );
  oai21d1 U2447 ( .B1(n1932), .B2(n1931), .A(n2290), .ZN(n3289) );
  inv0d0 U2448 ( .I(\hkspi/ldata[1] ), .ZN(n1934) );
  nr02d0 U2449 ( .A1(n2305), .A2(n2178), .ZN(n2179) );
  inv0d0 U2450 ( .I(n2179), .ZN(n2294) );
  oai222d1 U2451 ( .A1(n3289), .A2(n2298), .B1(n1934), .B2(n2296), .C1(n1933), 
        .C2(n2294), .ZN(n2547) );
  aoi22d1 U2452 ( .A1(n2282), .A2(\gpio_configure[9][10] ), .B1(n2238), .B2(
        \gpio_configure[3][10] ), .ZN(n1948) );
  aoi22d1 U2453 ( .A1(idata[0]), .A2(n2268), .B1(n2236), .B2(
        \gpio_configure[14][10] ), .ZN(n1947) );
  aoi22d1 U2454 ( .A1(n2252), .A2(\gpio_configure[37][10] ), .B1(n2230), .B2(
        \gpio_configure[4][10] ), .ZN(n1946) );
  aoi22d1 U2455 ( .A1(n2237), .A2(\gpio_configure[10][10] ), .B1(n2241), .B2(
        \gpio_configure[7][10] ), .ZN(n1938) );
  aoi22d1 U2456 ( .A1(n2257), .A2(\gpio_configure[35][10] ), .B1(n2224), .B2(
        \gpio_configure[12][10] ), .ZN(n1937) );
  aoi22d1 U2457 ( .A1(n2206), .A2(\gpio_configure[11][10] ), .B1(n2223), .B2(
        \gpio_configure[16][10] ), .ZN(n1936) );
  aoi22d1 U2458 ( .A1(n2231), .A2(\gpio_configure[34][10] ), .B1(n2222), .B2(
        \gpio_configure[5][10] ), .ZN(n1935) );
  aoi22d1 U2459 ( .A1(n2094), .A2(\gpio_configure[36][10] ), .B1(n2240), .B2(
        \gpio_configure[13][10] ), .ZN(n1942) );
  aoi22d1 U2460 ( .A1(n2242), .A2(\gpio_configure[2][10] ), .B1(n858), .B2(
        \gpio_configure[6][10] ), .ZN(n1941) );
  aoi22d1 U2461 ( .A1(n2251), .A2(mgmt_gpio_in[34]), .B1(n2281), .B2(
        \gpio_configure[8][10] ), .ZN(n1940) );
  aoi22d1 U2462 ( .A1(n2256), .A2(\gpio_configure[17][10] ), .B1(n844), .B2(
        \gpio_configure[15][10] ), .ZN(n1939) );
  nr02d0 U2463 ( .A1(n1944), .A2(n1943), .ZN(n1945) );
  aoi22d1 U2464 ( .A1(n2255), .A2(\gpio_configure[25][2] ), .B1(n2263), .B2(
        \gpio_configure[26][2] ), .ZN(n1951) );
  aoi22d1 U2465 ( .A1(n2253), .A2(\gpio_configure[27][2] ), .B1(n2225), .B2(
        \gpio_configure[19][2] ), .ZN(n1950) );
  aoi22d1 U2466 ( .A1(n2252), .A2(\gpio_configure[20][2] ), .B1(n2265), .B2(
        \gpio_configure[28][2] ), .ZN(n1949) );
  aoi211d1 U2467 ( .C1(n3229), .C2(pll_trim[10]), .A(n1953), .B(n1952), .ZN(
        n1997) );
  aoi22d1 U2468 ( .A1(n2206), .A2(pll_div[2]), .B1(n2041), .B2(
        \gpio_configure[18][2] ), .ZN(n1954) );
  oai21d1 U2469 ( .B1(n1956), .B2(n1955), .A(n1954), .ZN(n1962) );
  aoi22d1 U2470 ( .A1(n2276), .A2(\gpio_configure[31][2] ), .B1(n2200), .B2(
        \gpio_configure[22][2] ), .ZN(n1960) );
  aoi22d1 U2471 ( .A1(n2266), .A2(\gpio_configure[29][2] ), .B1(n2195), .B2(
        \gpio_configure[23][2] ), .ZN(n1959) );
  aoi22d1 U2472 ( .A1(n2254), .A2(\gpio_configure[32][2] ), .B1(n2001), .B2(
        \gpio_configure[21][2] ), .ZN(n1958) );
  aoi22d1 U2473 ( .A1(n2231), .A2(\gpio_configure[17][2] ), .B1(n2264), .B2(
        \gpio_configure[24][2] ), .ZN(n1957) );
  aoi211d1 U2474 ( .C1(n2256), .C2(\gpio_configure[0][2] ), .A(n1962), .B(
        n1961), .ZN(n1996) );
  aoi22d1 U2475 ( .A1(n2281), .A2(pll_trim[2]), .B1(n2258), .B2(
        \gpio_configure[31][10] ), .ZN(n1966) );
  aoi22d1 U2476 ( .A1(n2266), .A2(\gpio_configure[30][10] ), .B1(n2237), .B2(
        pll_sel[2]), .ZN(n1965) );
  aoi22d1 U2477 ( .A1(n2094), .A2(\gpio_configure[20][10] ), .B1(n2263), .B2(
        \gpio_configure[27][10] ), .ZN(n1964) );
  aoi22d1 U2478 ( .A1(n2268), .A2(\gpio_configure[24][10] ), .B1(n2257), .B2(
        \gpio_configure[19][10] ), .ZN(n1963) );
  aoi21d1 U2479 ( .B1(n2223), .B2(\gpio_configure[0][10] ), .A(n2242), .ZN(
        n1970) );
  aoi22d1 U2480 ( .A1(n2255), .A2(\gpio_configure[26][10] ), .B1(n844), .B2(
        clk1_output_dest), .ZN(n1969) );
  aoi22d1 U2481 ( .A1(n2269), .A2(\gpio_configure[23][10] ), .B1(n2264), .B2(
        \gpio_configure[25][10] ), .ZN(n1968) );
  aoi22d1 U2482 ( .A1(n2251), .A2(\gpio_configure[22][10] ), .B1(n2253), .B2(
        \gpio_configure[28][10] ), .ZN(n1967) );
  aoi22d1 U2483 ( .A1(n2282), .A2(pll_trim[18]), .B1(n2276), .B2(
        \gpio_configure[32][10] ), .ZN(n1974) );
  aoi22d1 U2484 ( .A1(n2256), .A2(\gpio_configure[1][10] ), .B1(n2252), .B2(
        \gpio_configure[21][10] ), .ZN(n1973) );
  aoi22d1 U2485 ( .A1(n2254), .A2(\gpio_configure[33][10] ), .B1(n2142), .B2(
        serial_bb_resetn), .ZN(n1972) );
  aoi22d1 U2486 ( .A1(n2265), .A2(\gpio_configure[29][10] ), .B1(n2267), .B2(
        \gpio_configure[18][10] ), .ZN(n1971) );
  aoim31d1 U2487 ( .B1(n1977), .B2(n1976), .B3(n1975), .A(n2288), .ZN(n1994)
         );
  aoi22d1 U2488 ( .A1(n2237), .A2(\gpio_configure[9][2] ), .B1(n2257), .B2(
        \gpio_configure[34][2] ), .ZN(n1981) );
  aoi22d1 U2489 ( .A1(n2223), .A2(\gpio_configure[15][2] ), .B1(n2240), .B2(
        \gpio_configure[12][2] ), .ZN(n1980) );
  aoi22d1 U2490 ( .A1(n2269), .A2(mgmt_gpio_in[26]), .B1(n2224), .B2(
        \gpio_configure[11][2] ), .ZN(n1979) );
  aoi22d1 U2491 ( .A1(n2264), .A2(n430), .B1(n2222), .B2(
        \gpio_configure[4][2] ), .ZN(n1978) );
  aoi22d1 U2492 ( .A1(n2252), .A2(\gpio_configure[36][2] ), .B1(n2242), .B2(
        \gpio_configure[1][2] ), .ZN(n1985) );
  aoi22d1 U2493 ( .A1(n2231), .A2(\gpio_configure[33][2] ), .B1(n2094), .B2(
        \gpio_configure[35][2] ), .ZN(n1984) );
  aoi22d1 U2494 ( .A1(n858), .A2(\gpio_configure[5][2] ), .B1(n2230), .B2(
        \gpio_configure[3][2] ), .ZN(n1983) );
  aoi22d1 U2495 ( .A1(n2256), .A2(\gpio_configure[16][2] ), .B1(n2236), .B2(
        \gpio_configure[13][2] ), .ZN(n1982) );
  aoi22d1 U2496 ( .A1(n3229), .A2(\gpio_configure[8][2] ), .B1(n844), .B2(
        \gpio_configure[14][2] ), .ZN(n1989) );
  aoi22d1 U2497 ( .A1(n2206), .A2(\gpio_configure[10][2] ), .B1(n2241), .B2(
        \gpio_configure[6][2] ), .ZN(n1988) );
  aoi22d1 U2498 ( .A1(n2251), .A2(\gpio_configure[37][2] ), .B1(n2281), .B2(
        \gpio_configure[7][2] ), .ZN(n1987) );
  aoi22d1 U2499 ( .A1(n2195), .A2(mgmt_gpio_in[10]), .B1(n2238), .B2(
        \gpio_configure[2][2] ), .ZN(n1986) );
  aoim31d1 U2500 ( .B1(n1992), .B2(n1991), .B3(n1990), .A(n2247), .ZN(n1993)
         );
  aoi211d1 U2501 ( .C1(n2283), .C2(mgmt_gpio_in[18]), .A(n1994), .B(n1993), 
        .ZN(n1995) );
  aon211d1 U2502 ( .C1(n1997), .C2(n1996), .B(n2277), .A(n1995), .ZN(n1998) );
  aon211d1 U2503 ( .C1(n2131), .C2(n1999), .B(n1998), .A(n2290), .ZN(n3285) );
  aoi22d1 U2504 ( .A1(\hkspi/ldata[1] ), .A2(n2179), .B1(\hkspi/ldata[2] ), 
        .B2(n2178), .ZN(n2000) );
  oai21d1 U2505 ( .B1(n3285), .B2(n2298), .A(n2000), .ZN(n2546) );
  aoi22d1 U2506 ( .A1(n2252), .A2(\gpio_configure[36][3] ), .B1(n2142), .B2(
        \gpio_configure[10][3] ), .ZN(n2015) );
  aoi22d1 U2507 ( .A1(n2267), .A2(\gpio_configure[33][3] ), .B1(n2001), .B2(
        \gpio_configure[37][3] ), .ZN(n2014) );
  aoi22d1 U2508 ( .A1(n2282), .A2(\gpio_configure[8][3] ), .B1(n2264), .B2(
        n429), .ZN(n2013) );
  aoi22d1 U2509 ( .A1(n2236), .A2(\gpio_configure[13][3] ), .B1(n2241), .B2(
        \gpio_configure[6][3] ), .ZN(n2005) );
  aoi22d1 U2510 ( .A1(n2094), .A2(\gpio_configure[35][3] ), .B1(n2224), .B2(
        \gpio_configure[11][3] ), .ZN(n2004) );
  aoi22d1 U2511 ( .A1(n2242), .A2(\gpio_configure[1][3] ), .B1(n2223), .B2(
        \gpio_configure[15][3] ), .ZN(n2003) );
  aoi22d1 U2512 ( .A1(n2256), .A2(\gpio_configure[16][3] ), .B1(n2238), .B2(
        \gpio_configure[2][3] ), .ZN(n2002) );
  aoi22d1 U2513 ( .A1(n858), .A2(\gpio_configure[5][3] ), .B1(n2230), .B2(
        \gpio_configure[3][3] ), .ZN(n2009) );
  aoi22d1 U2514 ( .A1(n2237), .A2(\gpio_configure[9][3] ), .B1(n2041), .B2(
        \gpio_configure[34][3] ), .ZN(n2008) );
  aoi22d1 U2515 ( .A1(n844), .A2(\gpio_configure[14][3] ), .B1(n2281), .B2(
        \gpio_configure[7][3] ), .ZN(n2007) );
  aoi22d1 U2516 ( .A1(n2240), .A2(\gpio_configure[12][3] ), .B1(n2222), .B2(
        \gpio_configure[4][3] ), .ZN(n2006) );
  nr02d0 U2517 ( .A1(n2011), .A2(n2010), .ZN(n2012) );
  aoi22d1 U2518 ( .A1(n2265), .A2(\gpio_configure[29][11] ), .B1(n2094), .B2(
        \gpio_configure[20][11] ), .ZN(n2018) );
  aoi22d1 U2519 ( .A1(n2282), .A2(pll_trim[19]), .B1(n2195), .B2(
        \gpio_configure[24][11] ), .ZN(n2017) );
  aoi22d1 U2520 ( .A1(n2251), .A2(\gpio_configure[22][11] ), .B1(n2266), .B2(
        \gpio_configure[30][11] ), .ZN(n2016) );
  aoi22d1 U2521 ( .A1(n2231), .A2(\gpio_configure[18][11] ), .B1(n2253), .B2(
        \gpio_configure[28][11] ), .ZN(n2022) );
  aoi22d1 U2522 ( .A1(n2256), .A2(\gpio_configure[1][11] ), .B1(n2263), .B2(
        \gpio_configure[27][11] ), .ZN(n2021) );
  aoi22d1 U2523 ( .A1(n2223), .A2(\gpio_configure[0][11] ), .B1(n2269), .B2(
        \gpio_configure[23][11] ), .ZN(n2020) );
  aoi22d1 U2524 ( .A1(n2255), .A2(\gpio_configure[26][11] ), .B1(n2237), .B2(
        pll90_sel[0]), .ZN(n2019) );
  aoi22d1 U2525 ( .A1(n2252), .A2(\gpio_configure[21][11] ), .B1(n2281), .B2(
        pll_trim[3]), .ZN(n2026) );
  aoi22d1 U2526 ( .A1(n2276), .A2(\gpio_configure[32][11] ), .B1(n2258), .B2(
        \gpio_configure[31][11] ), .ZN(n2025) );
  aoi22d1 U2527 ( .A1(n2254), .A2(\gpio_configure[33][11] ), .B1(n2264), .B2(
        \gpio_configure[25][11] ), .ZN(n2024) );
  aoi22d1 U2528 ( .A1(n2206), .A2(serial_bb_load), .B1(n2041), .B2(
        \gpio_configure[19][11] ), .ZN(n2023) );
  aoi22d1 U2529 ( .A1(n2285), .A2(mgmt_gpio_in[27]), .B1(n620), .B2(
        mgmt_gpio_in[11]), .ZN(n2062) );
  aoi22d1 U2530 ( .A1(n2258), .A2(\gpio_configure[30][3] ), .B1(n2094), .B2(
        \gpio_configure[19][3] ), .ZN(n2036) );
  aoi22d1 U2531 ( .A1(n2256), .A2(\gpio_configure[0][3] ), .B1(n2253), .B2(
        \gpio_configure[27][3] ), .ZN(n2035) );
  aoi22d1 U2532 ( .A1(n2265), .A2(\gpio_configure[28][3] ), .B1(n2142), .B2(
        pll_div[3]), .ZN(n2032) );
  inv0d0 U2533 ( .I(n2076), .ZN(n2239) );
  aoi22d1 U2534 ( .A1(n2239), .A2(\gpio_configure[20][3] ), .B1(n2251), .B2(
        \gpio_configure[21][3] ), .ZN(n2031) );
  aoi22d1 U2535 ( .A1(n2266), .A2(\gpio_configure[29][3] ), .B1(n2195), .B2(
        \gpio_configure[23][3] ), .ZN(n2030) );
  aoi211d1 U2536 ( .C1(n3229), .C2(pll_trim[11]), .A(n844), .B(n2033), .ZN(
        n2034) );
  aoi22d1 U2537 ( .A1(n2276), .A2(\gpio_configure[31][3] ), .B1(n2267), .B2(
        \gpio_configure[17][3] ), .ZN(n2040) );
  aoi22d1 U2538 ( .A1(n2254), .A2(\gpio_configure[32][3] ), .B1(n2269), .B2(
        \gpio_configure[22][3] ), .ZN(n2039) );
  aoi22d1 U2539 ( .A1(n2264), .A2(\gpio_configure[24][3] ), .B1(n2041), .B2(
        \gpio_configure[18][3] ), .ZN(n2038) );
  aoi22d1 U2540 ( .A1(n2255), .A2(\gpio_configure[25][3] ), .B1(n2263), .B2(
        \gpio_configure[26][3] ), .ZN(n2037) );
  aoi22d1 U2541 ( .A1(n2206), .A2(\gpio_configure[11][11] ), .B1(n2041), .B2(
        \gpio_configure[35][11] ), .ZN(n2057) );
  aoi22d1 U2542 ( .A1(n2269), .A2(mgmt_gpio_in[19]), .B1(n2222), .B2(
        \gpio_configure[5][11] ), .ZN(n2056) );
  aoi22d1 U2543 ( .A1(n858), .A2(\gpio_configure[6][11] ), .B1(n2230), .B2(
        \gpio_configure[4][11] ), .ZN(n2053) );
  aoi22d1 U2544 ( .A1(n2223), .A2(\gpio_configure[16][11] ), .B1(n844), .B2(
        \gpio_configure[15][11] ), .ZN(n2052) );
  aoi22d1 U2545 ( .A1(n2238), .A2(\gpio_configure[3][11] ), .B1(n2241), .B2(
        \gpio_configure[7][11] ), .ZN(n2044) );
  aoi22d1 U2546 ( .A1(n2282), .A2(\gpio_configure[9][11] ), .B1(n2240), .B2(
        \gpio_configure[13][11] ), .ZN(n2043) );
  aoi22d1 U2547 ( .A1(n2251), .A2(mgmt_gpio_in[35]), .B1(n2236), .B2(
        \gpio_configure[14][11] ), .ZN(n2042) );
  aoi22d1 U2548 ( .A1(n2256), .A2(\gpio_configure[17][11] ), .B1(n2224), .B2(
        \gpio_configure[12][11] ), .ZN(n2048) );
  aoi22d1 U2549 ( .A1(n2237), .A2(\gpio_configure[10][11] ), .B1(n2094), .B2(
        \gpio_configure[36][11] ), .ZN(n2047) );
  aoi22d1 U2550 ( .A1(n2242), .A2(\gpio_configure[2][11] ), .B1(n2281), .B2(
        \gpio_configure[8][11] ), .ZN(n2046) );
  aoi22d1 U2551 ( .A1(n2239), .A2(\gpio_configure[37][11] ), .B1(n2195), .B2(
        mgmt_gpio_in[3]), .ZN(n2045) );
  aoi211d1 U2552 ( .C1(n2267), .C2(\gpio_configure[34][11] ), .A(n2050), .B(
        n2049), .ZN(n2051) );
  an03d0 U2553 ( .A1(n2053), .A2(n2052), .A3(n2051), .Z(n2055) );
  aoi31d1 U2554 ( .B1(n2057), .B2(n2056), .B3(n2055), .A(n2054), .ZN(n2058) );
  oan211d1 U2555 ( .C1(n2060), .C2(n2059), .B(n2220), .A(n2058), .ZN(n2061) );
  oai211d1 U2556 ( .C1(n2063), .C2(n2288), .A(n2062), .B(n2061), .ZN(n2064) );
  aon211d1 U2557 ( .C1(n2211), .C2(n2065), .B(n2064), .A(n2290), .ZN(n3284) );
  aoi22d1 U2558 ( .A1(\hkspi/ldata[2] ), .A2(n2179), .B1(\hkspi/ldata[3] ), 
        .B2(n2178), .ZN(n2066) );
  oai21d1 U2559 ( .B1(n2298), .B2(n3284), .A(n2066), .ZN(n2545) );
  aoi22d1 U2560 ( .A1(n2068), .A2(\gpio_configure[0][12] ), .B1(n2067), .B2(
        pll90_sel[1]), .ZN(n2086) );
  aoi22d1 U2561 ( .A1(n2256), .A2(\gpio_configure[1][12] ), .B1(n2263), .B2(
        \gpio_configure[27][12] ), .ZN(n2085) );
  aoi22d1 U2562 ( .A1(n2231), .A2(\gpio_configure[18][12] ), .B1(n2255), .B2(
        \gpio_configure[26][12] ), .ZN(n2070) );
  aoi22d1 U2563 ( .A1(n2251), .A2(\gpio_configure[22][12] ), .B1(n2258), .B2(
        \gpio_configure[31][12] ), .ZN(n2069) );
  oai211d1 U2564 ( .C1(n2072), .C2(n2071), .A(n2070), .B(n2069), .ZN(n2073) );
  aoi211d1 U2565 ( .C1(n2195), .C2(\gpio_configure[24][12] ), .A(n2238), .B(
        n2073), .ZN(n2084) );
  aoi22d1 U2566 ( .A1(n2254), .A2(\gpio_configure[33][12] ), .B1(n2281), .B2(
        pll_trim[4]), .ZN(n2074) );
  oai21d1 U2567 ( .B1(n2076), .B2(n2075), .A(n2074), .ZN(n2082) );
  aoi22d1 U2568 ( .A1(n2269), .A2(\gpio_configure[23][12] ), .B1(n2264), .B2(
        \gpio_configure[25][12] ), .ZN(n2080) );
  aoi22d1 U2569 ( .A1(n3229), .A2(pll_trim[20]), .B1(n2266), .B2(
        \gpio_configure[30][12] ), .ZN(n2079) );
  aoi22d1 U2570 ( .A1(n2276), .A2(\gpio_configure[32][12] ), .B1(n2094), .B2(
        \gpio_configure[20][12] ), .ZN(n2078) );
  aoi22d1 U2571 ( .A1(n2206), .A2(serial_bb_clock), .B1(n2253), .B2(
        \gpio_configure[28][12] ), .ZN(n2077) );
  aoi211d1 U2572 ( .C1(n2265), .C2(\gpio_configure[29][12] ), .A(n2082), .B(
        n2081), .ZN(n2083) );
  aoi22d1 U2573 ( .A1(n2206), .A2(pll_div[4]), .B1(n2266), .B2(
        \gpio_configure[29][4] ), .ZN(n2089) );
  aoi22d1 U2574 ( .A1(n2282), .A2(pll_trim[12]), .B1(n2251), .B2(
        \gpio_configure[21][4] ), .ZN(n2088) );
  aoi22d1 U2575 ( .A1(n2265), .A2(\gpio_configure[28][4] ), .B1(n2255), .B2(
        \gpio_configure[25][4] ), .ZN(n2087) );
  aoi211d1 U2576 ( .C1(n2263), .C2(\gpio_configure[26][4] ), .A(n2238), .B(
        n2090), .ZN(n2134) );
  aoi22d1 U2577 ( .A1(n2254), .A2(\gpio_configure[32][4] ), .B1(n2258), .B2(
        \gpio_configure[30][4] ), .ZN(n2091) );
  oai21d1 U2578 ( .B1(n2093), .B2(n2092), .A(n2091), .ZN(n2100) );
  aoi22d1 U2579 ( .A1(n2239), .A2(\gpio_configure[20][4] ), .B1(n2200), .B2(
        \gpio_configure[22][4] ), .ZN(n2098) );
  aoi22d1 U2580 ( .A1(n2276), .A2(\gpio_configure[31][4] ), .B1(n2264), .B2(
        \gpio_configure[24][4] ), .ZN(n2097) );
  aoi22d1 U2581 ( .A1(n2253), .A2(\gpio_configure[27][4] ), .B1(n2257), .B2(
        \gpio_configure[18][4] ), .ZN(n2096) );
  aoi22d1 U2582 ( .A1(n2231), .A2(\gpio_configure[17][4] ), .B1(n2094), .B2(
        \gpio_configure[19][4] ), .ZN(n2095) );
  aoi211d1 U2583 ( .C1(n2256), .C2(\gpio_configure[0][4] ), .A(n2100), .B(
        n2099), .ZN(n2133) );
  aoi22d1 U2584 ( .A1(n3229), .A2(\gpio_configure[9][12] ), .B1(n2240), .B2(
        \gpio_configure[13][12] ), .ZN(n2114) );
  aoi22d1 U2585 ( .A1(n844), .A2(\gpio_configure[15][12] ), .B1(n2236), .B2(
        \gpio_configure[14][12] ), .ZN(n2113) );
  aoi22d1 U2586 ( .A1(n2225), .A2(\gpio_configure[36][12] ), .B1(n2238), .B2(
        \gpio_configure[3][12] ), .ZN(n2112) );
  aoi22d1 U2587 ( .A1(n2239), .A2(\gpio_configure[37][12] ), .B1(n2230), .B2(
        \gpio_configure[4][12] ), .ZN(n2104) );
  aoi22d1 U2588 ( .A1(n2256), .A2(\gpio_configure[17][12] ), .B1(n2237), .B2(
        \gpio_configure[10][12] ), .ZN(n2103) );
  aoi22d1 U2589 ( .A1(n2231), .A2(\gpio_configure[34][12] ), .B1(n2224), .B2(
        \gpio_configure[12][12] ), .ZN(n2102) );
  aoi22d1 U2590 ( .A1(n858), .A2(\gpio_configure[6][12] ), .B1(n2241), .B2(
        \gpio_configure[7][12] ), .ZN(n2101) );
  aoi22d1 U2591 ( .A1(n2269), .A2(mgmt_gpio_in[20]), .B1(n2257), .B2(
        \gpio_configure[35][12] ), .ZN(n2108) );
  aoi22d1 U2592 ( .A1(n2206), .A2(\gpio_configure[11][12] ), .B1(n2242), .B2(
        \gpio_configure[2][12] ), .ZN(n2107) );
  aoi22d1 U2593 ( .A1(n2281), .A2(\gpio_configure[8][12] ), .B1(n2222), .B2(
        \gpio_configure[5][12] ), .ZN(n2106) );
  aoi22d1 U2594 ( .A1(n2223), .A2(\gpio_configure[16][12] ), .B1(n2251), .B2(
        mgmt_gpio_in[36]), .ZN(n2105) );
  nr02d0 U2595 ( .A1(n2110), .A2(n2109), .ZN(n2111) );
  aoi22d1 U2596 ( .A1(n2239), .A2(\gpio_configure[36][4] ), .B1(n858), .B2(
        \gpio_configure[5][4] ), .ZN(n2118) );
  aoi22d1 U2597 ( .A1(n2242), .A2(\gpio_configure[1][4] ), .B1(n2223), .B2(
        \gpio_configure[15][4] ), .ZN(n2117) );
  aoi22d1 U2598 ( .A1(n2225), .A2(\gpio_configure[35][4] ), .B1(n2241), .B2(
        \gpio_configure[6][4] ), .ZN(n2116) );
  aoi22d1 U2599 ( .A1(n2238), .A2(\gpio_configure[2][4] ), .B1(n2224), .B2(
        \gpio_configure[11][4] ), .ZN(n2115) );
  aoi22d1 U2600 ( .A1(n2269), .A2(mgmt_gpio_in[28]), .B1(n2257), .B2(
        \gpio_configure[34][4] ), .ZN(n2121) );
  aoi22d1 U2601 ( .A1(n2256), .A2(\gpio_configure[16][4] ), .B1(n844), .B2(
        \gpio_configure[14][4] ), .ZN(n2120) );
  aoi22d1 U2602 ( .A1(n3229), .A2(\gpio_configure[8][4] ), .B1(n2240), .B2(
        \gpio_configure[12][4] ), .ZN(n2119) );
  aoi22d1 U2603 ( .A1(n2231), .A2(\gpio_configure[33][4] ), .B1(n2142), .B2(
        \gpio_configure[10][4] ), .ZN(n2125) );
  aoi22d1 U2604 ( .A1(n2251), .A2(\gpio_configure[37][4] ), .B1(n2222), .B2(
        \gpio_configure[4][4] ), .ZN(n2124) );
  aoi22d1 U2605 ( .A1(n2237), .A2(\gpio_configure[9][4] ), .B1(n2230), .B2(
        \gpio_configure[3][4] ), .ZN(n2123) );
  aoi22d1 U2606 ( .A1(n2281), .A2(\gpio_configure[7][4] ), .B1(n2236), .B2(
        \gpio_configure[13][4] ), .ZN(n2122) );
  aoim31d1 U2607 ( .B1(n2128), .B2(n2127), .B3(n2126), .A(n2247), .ZN(n2129)
         );
  aoi211d1 U2608 ( .C1(n2131), .C2(n2130), .A(n2129), .B(n386), .ZN(n2132) );
  aon211d1 U2609 ( .C1(n2134), .C2(n2133), .B(n2277), .A(n2132), .ZN(n2135) );
  aon211d1 U2610 ( .C1(n2137), .C2(n2136), .B(n2135), .A(n2290), .ZN(n3280) );
  aoi22d1 U2611 ( .A1(\hkspi/ldata[3] ), .A2(n2179), .B1(\hkspi/ldata[4] ), 
        .B2(n2178), .ZN(n2138) );
  oai21d1 U2612 ( .B1(n2298), .B2(n3280), .A(n2138), .ZN(n2544) );
  mx02d1 U2613 ( .I0(serial_bb_data_1), .I1(serial_data_staging_1[12]), .S(
        n2181), .Z(serial_data_1) );
  aoi22d1 U2614 ( .A1(n2285), .A2(mgmt_gpio_in[29]), .B1(n2139), .B2(
        mgmt_gpio_in[37]), .ZN(n2141) );
  aoi22d1 U2615 ( .A1(n2283), .A2(mgmt_gpio_in[21]), .B1(n620), .B2(
        mgmt_gpio_in[13]), .ZN(n2140) );
  oaim211d1 U2616 ( .C1(mgmt_gpio_in[5]), .C2(n2284), .A(n2141), .B(n2140), 
        .ZN(n2177) );
  aoi22d1 U2617 ( .A1(n3229), .A2(pll_trim[21]), .B1(n2142), .B2(serial_data_1), .ZN(n2160) );
  aoi22d1 U2618 ( .A1(n2281), .A2(pll_trim[5]), .B1(n2237), .B2(pll90_sel[2]), 
        .ZN(n2159) );
  aoi22d1 U2619 ( .A1(n2256), .A2(\gpio_configure[16][5] ), .B1(n2251), .B2(
        \gpio_configure[37][5] ), .ZN(n2146) );
  aoi22d1 U2620 ( .A1(n2206), .A2(\gpio_configure[10][5] ), .B1(n2242), .B2(
        \gpio_configure[1][5] ), .ZN(n2145) );
  aoi22d1 U2621 ( .A1(n2225), .A2(\gpio_configure[35][5] ), .B1(n2222), .B2(
        \gpio_configure[4][5] ), .ZN(n2144) );
  aoi22d1 U2622 ( .A1(n2223), .A2(\gpio_configure[15][5] ), .B1(n2224), .B2(
        \gpio_configure[11][5] ), .ZN(n2143) );
  aoi22d1 U2623 ( .A1(n2231), .A2(\gpio_configure[33][5] ), .B1(n2230), .B2(
        \gpio_configure[3][5] ), .ZN(n2148) );
  aoi22d1 U2624 ( .A1(n2281), .A2(\gpio_configure[7][5] ), .B1(n858), .B2(
        \gpio_configure[5][5] ), .ZN(n2147) );
  oai211d1 U2625 ( .C1(n2150), .C2(n2149), .A(n2148), .B(n2147), .ZN(n2156) );
  aoi22d1 U2626 ( .A1(n2237), .A2(\gpio_configure[9][5] ), .B1(n2236), .B2(
        \gpio_configure[13][5] ), .ZN(n2154) );
  aoi22d1 U2627 ( .A1(n2239), .A2(\gpio_configure[36][5] ), .B1(n844), .B2(
        \gpio_configure[14][5] ), .ZN(n2153) );
  aoi22d1 U2628 ( .A1(n2257), .A2(\gpio_configure[34][5] ), .B1(n2241), .B2(
        \gpio_configure[6][5] ), .ZN(n2152) );
  aoi22d1 U2629 ( .A1(n3229), .A2(\gpio_configure[8][5] ), .B1(n2240), .B2(
        \gpio_configure[12][5] ), .ZN(n2151) );
  oai31d1 U2630 ( .B1(n2157), .B2(n2156), .B3(n2155), .A(n2211), .ZN(n2158) );
  aon211d1 U2631 ( .C1(n2160), .C2(n2159), .B(n2288), .A(n2158), .ZN(n2176) );
  aoi22d1 U2632 ( .A1(n2254), .A2(\gpio_configure[32][5] ), .B1(n2255), .B2(
        \gpio_configure[25][5] ), .ZN(n2174) );
  aoi22d1 U2633 ( .A1(n2282), .A2(pll_trim[13]), .B1(n2253), .B2(
        \gpio_configure[27][5] ), .ZN(n2173) );
  aoi22d1 U2634 ( .A1(n2264), .A2(\gpio_configure[24][5] ), .B1(n2251), .B2(
        \gpio_configure[21][5] ), .ZN(n2162) );
  aoi22d1 U2635 ( .A1(n2225), .A2(\gpio_configure[19][5] ), .B1(n2195), .B2(
        \gpio_configure[23][5] ), .ZN(n2161) );
  oai211d1 U2636 ( .C1(n2164), .C2(n2163), .A(n2162), .B(n2161), .ZN(n2170) );
  aoi22d1 U2637 ( .A1(n2265), .A2(\gpio_configure[28][5] ), .B1(n2266), .B2(
        \gpio_configure[29][5] ), .ZN(n2168) );
  aoi22d1 U2638 ( .A1(n2239), .A2(\gpio_configure[20][5] ), .B1(n2258), .B2(
        \gpio_configure[30][5] ), .ZN(n2167) );
  aoi22d1 U2639 ( .A1(n2276), .A2(\gpio_configure[31][5] ), .B1(n2263), .B2(
        \gpio_configure[26][5] ), .ZN(n2166) );
  aoi22d1 U2640 ( .A1(n2269), .A2(\gpio_configure[22][5] ), .B1(n2257), .B2(
        \gpio_configure[18][5] ), .ZN(n2165) );
  aoi211d1 U2641 ( .C1(n2267), .C2(\gpio_configure[17][5] ), .A(n2170), .B(
        n2169), .ZN(n2172) );
  aoi31d1 U2642 ( .B1(n2174), .B2(n2173), .B3(n2172), .A(n2171), .ZN(n2175) );
  oan211d1 U2643 ( .C1(n2177), .C2(n2176), .B(n2290), .A(n2175), .ZN(n3281) );
  aoi22d1 U2644 ( .A1(\hkspi/ldata[4] ), .A2(n2179), .B1(\hkspi/ldata[5] ), 
        .B2(n2178), .ZN(n2180) );
  oai21d1 U2645 ( .B1(n3281), .B2(n2298), .A(n2180), .ZN(n2543) );
  mx02d1 U2646 ( .I0(serial_bb_data_2), .I1(serial_data_staging_2[12]), .S(
        n2181), .Z(serial_data_2) );
  inv0d0 U2647 ( .I(\hkspi/ldata[5] ), .ZN(n2221) );
  inv0d0 U2648 ( .I(\hkspi/ldata[6] ), .ZN(n2295) );
  aoi22d1 U2649 ( .A1(n2256), .A2(\gpio_configure[0][6] ), .B1(n2257), .B2(
        \gpio_configure[18][6] ), .ZN(n2194) );
  aoi22d1 U2650 ( .A1(n2254), .A2(\gpio_configure[32][6] ), .B1(n2258), .B2(
        \gpio_configure[30][6] ), .ZN(n2193) );
  aoi22d1 U2651 ( .A1(n2253), .A2(\gpio_configure[27][6] ), .B1(n2266), .B2(
        \gpio_configure[29][6] ), .ZN(n2183) );
  aoi22d1 U2652 ( .A1(n2225), .A2(\gpio_configure[19][6] ), .B1(n2195), .B2(
        \gpio_configure[23][6] ), .ZN(n2182) );
  oai211d1 U2653 ( .C1(n2185), .C2(n2184), .A(n2183), .B(n2182), .ZN(n2186) );
  aoi211d1 U2654 ( .C1(n2200), .C2(\gpio_configure[22][6] ), .A(n2238), .B(
        n2186), .ZN(n2192) );
  aoi22d1 U2655 ( .A1(n2239), .A2(\gpio_configure[20][6] ), .B1(n2276), .B2(
        \gpio_configure[31][6] ), .ZN(n2190) );
  aoi22d1 U2656 ( .A1(n2282), .A2(pll_trim[14]), .B1(n2263), .B2(
        \gpio_configure[26][6] ), .ZN(n2189) );
  aoi22d1 U2657 ( .A1(n2265), .A2(\gpio_configure[28][6] ), .B1(n2255), .B2(
        \gpio_configure[25][6] ), .ZN(n2188) );
  aoi22d1 U2658 ( .A1(n2231), .A2(\gpio_configure[17][6] ), .B1(n2251), .B2(
        \gpio_configure[21][6] ), .ZN(n2187) );
  an04d0 U2659 ( .A1(n2190), .A2(n2189), .A3(n2188), .A4(n2187), .Z(n2191) );
  aoi222d1 U2660 ( .A1(serial_data_2), .A2(n2206), .B1(n2281), .B2(pll_trim[6]), .C1(n2282), .C2(pll_trim[22]), .ZN(n2217) );
  aoi22d1 U2661 ( .A1(n2283), .A2(mgmt_gpio_in[22]), .B1(n2284), .B2(
        mgmt_gpio_in[6]), .ZN(n2216) );
  aoi22d1 U2662 ( .A1(n2256), .A2(\gpio_configure[16][6] ), .B1(n2252), .B2(
        \gpio_configure[36][6] ), .ZN(n2199) );
  aoi22d1 U2663 ( .A1(n2231), .A2(\gpio_configure[33][6] ), .B1(n2238), .B2(
        \gpio_configure[2][6] ), .ZN(n2198) );
  aoi22d1 U2664 ( .A1(n2195), .A2(mgmt_gpio_in[14]), .B1(n2240), .B2(
        \gpio_configure[12][6] ), .ZN(n2197) );
  aoi22d1 U2665 ( .A1(n2242), .A2(\gpio_configure[1][6] ), .B1(n844), .B2(
        \gpio_configure[14][6] ), .ZN(n2196) );
  aoi22d1 U2666 ( .A1(n2223), .A2(\gpio_configure[15][6] ), .B1(n2257), .B2(
        \gpio_configure[34][6] ), .ZN(n2204) );
  aoi22d1 U2667 ( .A1(n2282), .A2(\gpio_configure[8][6] ), .B1(n2224), .B2(
        \gpio_configure[11][6] ), .ZN(n2203) );
  aoi22d1 U2668 ( .A1(n2237), .A2(\gpio_configure[9][6] ), .B1(n858), .B2(
        \gpio_configure[5][6] ), .ZN(n2202) );
  nd02d0 U2669 ( .A1(n2200), .A2(mgmt_gpio_in[30]), .ZN(n2201) );
  aoi22d1 U2670 ( .A1(n2205), .A2(\gpio_configure[7][6] ), .B1(n2241), .B2(
        \gpio_configure[6][6] ), .ZN(n2210) );
  aoi22d1 U2671 ( .A1(n2225), .A2(\gpio_configure[35][6] ), .B1(n2236), .B2(
        \gpio_configure[13][6] ), .ZN(n2209) );
  aoi22d1 U2672 ( .A1(n2206), .A2(\gpio_configure[10][6] ), .B1(n2222), .B2(
        \gpio_configure[4][6] ), .ZN(n2208) );
  aoi22d1 U2673 ( .A1(n2251), .A2(\gpio_configure[37][6] ), .B1(n2230), .B2(
        \gpio_configure[3][6] ), .ZN(n2207) );
  oai31d1 U2674 ( .B1(n2214), .B2(n2213), .B3(n2212), .A(n2211), .ZN(n2215) );
  oai211d1 U2675 ( .C1(n2217), .C2(n2288), .A(n2216), .B(n2215), .ZN(n2218) );
  aon211d1 U2676 ( .C1(n2220), .C2(n2219), .B(n2218), .A(n2290), .ZN(n3282) );
  oai222d1 U2677 ( .A1(n2294), .A2(n2221), .B1(n2295), .B2(n2296), .C1(n2298), 
        .C2(n3282), .ZN(n2542) );
  aoi22d1 U2678 ( .A1(n2282), .A2(\gpio_configure[8][7] ), .B1(n2251), .B2(
        \gpio_configure[37][7] ), .ZN(n2229) );
  aoi22d1 U2679 ( .A1(n2223), .A2(\gpio_configure[15][7] ), .B1(n2222), .B2(
        \gpio_configure[4][7] ), .ZN(n2228) );
  aoi22d1 U2680 ( .A1(n2256), .A2(\gpio_configure[16][7] ), .B1(n2224), .B2(
        \gpio_configure[11][7] ), .ZN(n2227) );
  aoi22d1 U2681 ( .A1(n2225), .A2(\gpio_configure[35][7] ), .B1(n858), .B2(
        \gpio_configure[5][7] ), .ZN(n2226) );
  aoi22d1 U2682 ( .A1(n844), .A2(\gpio_configure[14][7] ), .B1(n2230), .B2(
        \gpio_configure[3][7] ), .ZN(n2233) );
  aoi22d1 U2683 ( .A1(n2231), .A2(\gpio_configure[33][7] ), .B1(n2257), .B2(
        \gpio_configure[34][7] ), .ZN(n2232) );
  oai211d1 U2684 ( .C1(n2235), .C2(n2234), .A(n2233), .B(n2232), .ZN(n2249) );
  aoi22d1 U2685 ( .A1(n2237), .A2(\gpio_configure[9][7] ), .B1(n2236), .B2(
        \gpio_configure[13][7] ), .ZN(n2246) );
  aoi22d1 U2686 ( .A1(n2239), .A2(\gpio_configure[36][7] ), .B1(n2238), .B2(
        \gpio_configure[2][7] ), .ZN(n2245) );
  aoi22d1 U2687 ( .A1(n2281), .A2(\gpio_configure[7][7] ), .B1(n2240), .B2(
        \gpio_configure[12][7] ), .ZN(n2244) );
  aoi22d1 U2688 ( .A1(n2242), .A2(\gpio_configure[1][7] ), .B1(n2241), .B2(
        \gpio_configure[6][7] ), .ZN(n2243) );
  aoim31d1 U2689 ( .B1(n2250), .B2(n2249), .B3(n2248), .A(n2247), .ZN(n2293)
         );
  aoi22d1 U2690 ( .A1(n2252), .A2(\gpio_configure[20][7] ), .B1(n2251), .B2(
        \gpio_configure[21][7] ), .ZN(n2280) );
  aoi22d1 U2691 ( .A1(n2254), .A2(\gpio_configure[32][7] ), .B1(n2253), .B2(
        \gpio_configure[27][7] ), .ZN(n2279) );
  aoi22d1 U2692 ( .A1(n2256), .A2(\gpio_configure[0][7] ), .B1(n2255), .B2(
        \gpio_configure[25][7] ), .ZN(n2260) );
  aoi22d1 U2693 ( .A1(n2258), .A2(\gpio_configure[30][7] ), .B1(n2257), .B2(
        \gpio_configure[18][7] ), .ZN(n2259) );
  oai211d1 U2694 ( .C1(n2262), .C2(n2261), .A(n2260), .B(n2259), .ZN(n2275) );
  aoi22d1 U2695 ( .A1(n2264), .A2(\gpio_configure[24][7] ), .B1(n2263), .B2(
        \gpio_configure[26][7] ), .ZN(n2273) );
  aoi22d1 U2696 ( .A1(n3229), .A2(pll_trim[15]), .B1(n2265), .B2(
        \gpio_configure[28][7] ), .ZN(n2272) );
  aoi22d1 U2697 ( .A1(n2267), .A2(\gpio_configure[17][7] ), .B1(n2266), .B2(
        \gpio_configure[29][7] ), .ZN(n2271) );
  aoi22d1 U2698 ( .A1(n2269), .A2(\gpio_configure[22][7] ), .B1(n2268), .B2(
        \gpio_configure[23][7] ), .ZN(n2270) );
  aoi211d1 U2699 ( .C1(n2276), .C2(\gpio_configure[31][7] ), .A(n2275), .B(
        n2274), .ZN(n2278) );
  aoi31d1 U2700 ( .B1(n2280), .B2(n2279), .B3(n2278), .A(n2277), .ZN(n2292) );
  aoi22d1 U2701 ( .A1(n2282), .A2(pll_trim[23]), .B1(n2281), .B2(pll_trim[7]), 
        .ZN(n2289) );
  aoi22d1 U2702 ( .A1(n2283), .A2(mgmt_gpio_in[23]), .B1(n620), .B2(
        mgmt_gpio_in[15]), .ZN(n2287) );
  aoi22d1 U2703 ( .A1(n2285), .A2(mgmt_gpio_in[31]), .B1(n2284), .B2(
        mgmt_gpio_in[7]), .ZN(n2286) );
  oai211d1 U2704 ( .C1(n2289), .C2(n2288), .A(n2287), .B(n2286), .ZN(n2291) );
  oai31d1 U2705 ( .B1(n2293), .B2(n2292), .B3(n2291), .A(n2290), .ZN(n3279) );
  oai222d1 U2706 ( .A1(n3279), .A2(n2298), .B1(n2297), .B2(n2296), .C1(n2295), 
        .C2(n2294), .ZN(n2541) );
  aoim22d1 U2708 ( .A1(n2302), .A2(n2301), .B1(n2300), .B2(n2299), .Z(n2534)
         );
  aoim22d1 U2709 ( .A1(n2304), .A2(n2303), .B1(n2303), .B2(
        \hkspi/pre_pass_thru_user ), .Z(n2533) );
  nd12d0 U2710 ( .A1(n2316), .A2(n2305), .ZN(n2306) );
  mx02d1 U2711 ( .I0(idata[0]), .I1(\hkspi/writemode ), .S(n2306), .Z(n2532)
         );
  inv0d0 U2712 ( .I(idata[1]), .ZN(n2308) );
  aoi22d1 U2713 ( .A1(n2315), .A2(n2307), .B1(n2308), .B2(n2312), .ZN(n2531)
         );
  inv0d0 U2714 ( .I(idata[2]), .ZN(n2309) );
  aoi22d1 U2715 ( .A1(n2315), .A2(n2308), .B1(n2309), .B2(n2312), .ZN(n2530)
         );
  inv0d0 U2716 ( .I(idata[3]), .ZN(n2310) );
  aoi22d1 U2717 ( .A1(n2315), .A2(n2309), .B1(n2310), .B2(n2312), .ZN(n2529)
         );
  inv0d0 U2718 ( .I(idata[4]), .ZN(n2311) );
  aoi22d1 U2719 ( .A1(n2315), .A2(n2310), .B1(n2311), .B2(n2312), .ZN(n2528)
         );
  inv0d0 U2720 ( .I(idata[5]), .ZN(n2313) );
  aoi22d1 U2721 ( .A1(n2315), .A2(n2311), .B1(n2313), .B2(n2312), .ZN(n2527)
         );
  inv0d0 U2722 ( .I(idata[6]), .ZN(n2314) );
  aoi22d1 U2723 ( .A1(n2315), .A2(n2313), .B1(n2314), .B2(n2312), .ZN(n2526)
         );
  aoim22d1 U2724 ( .A1(n2315), .A2(n2314), .B1(idata[7]), .B2(n2315), .Z(n2525) );
  nr04d0 U2725 ( .A1(\hkspi/count[2] ), .A2(\hkspi/count[1] ), .A3(n2317), 
        .A4(n2316), .ZN(n2318) );
  mx02d1 U2726 ( .I0(\hkspi/readmode ), .I1(idata[0]), .S(n2318), .Z(n2524) );
  inv0d0 U2727 ( .I(n2321), .ZN(n2320) );
  aoi22d1 U2728 ( .A1(n2321), .A2(n3157), .B1(\gpio_configure[4][10] ), .B2(
        n2320), .ZN(n2522) );
  inv0d0 U2729 ( .I(n2324), .ZN(n2323) );
  aoi22d1 U2730 ( .A1(n2324), .A2(n3157), .B1(\gpio_configure[16][10] ), .B2(
        n2323), .ZN(n2521) );
  inv0d0 U2731 ( .I(n2326), .ZN(n2325) );
  aoi22d1 U2732 ( .A1(n2326), .A2(n3242), .B1(\gpio_configure[15][1] ), .B2(
        n2325), .ZN(n2520) );
  aoi22d1 U2733 ( .A1(n2326), .A2(n3233), .B1(\gpio_configure[15][0] ), .B2(
        n2325), .ZN(n2519) );
  aoi22d1 U2734 ( .A1(n2328), .A2(n3230), .B1(\gpio_configure[0][12] ), .B2(
        n2327), .ZN(n2518) );
  aoi22d1 U2735 ( .A1(n2328), .A2(n3231), .B1(\gpio_configure[0][11] ), .B2(
        n2327), .ZN(n2517) );
  aoi22d1 U2736 ( .A1(n2330), .A2(n3157), .B1(\gpio_configure[8][10] ), .B2(
        n2329), .ZN(n2516) );
  inv0d0 U2737 ( .I(n2332), .ZN(n2331) );
  aoi22d1 U2738 ( .A1(n2332), .A2(n3242), .B1(\gpio_configure[7][1] ), .B2(
        n2331), .ZN(n2515) );
  aoi22d1 U2739 ( .A1(n2332), .A2(n3233), .B1(\gpio_configure[7][0] ), .B2(
        n2331), .ZN(n2514) );
  nr02d0 U2740 ( .A1(n2334), .A2(n2333), .ZN(n2337) );
  inv0d0 U2741 ( .I(n2337), .ZN(n2336) );
  aoi22d1 U2742 ( .A1(n2336), .A2(pll_trim[7]), .B1(n3235), .B2(n2337), .ZN(
        n2513) );
  aoi22d1 U2743 ( .A1(n2337), .A2(n3236), .B1(pll_trim[6]), .B2(n2336), .ZN(
        n2512) );
  aoi22d1 U2744 ( .A1(n2337), .A2(n3237), .B1(pll_trim[5]), .B2(n2336), .ZN(
        n2511) );
  aoi22d1 U2745 ( .A1(n2337), .A2(n3230), .B1(pll_trim[4]), .B2(n2336), .ZN(
        n2510) );
  aoi22d1 U2746 ( .A1(n2337), .A2(n3231), .B1(pll_trim[3]), .B2(n2336), .ZN(
        n2509) );
  aoi22d1 U2747 ( .A1(n2337), .A2(n3157), .B1(pll_trim[2]), .B2(n2336), .ZN(
        n2508) );
  aoi22d1 U2748 ( .A1(n2337), .A2(n3242), .B1(pll_trim[1]), .B2(n2336), .ZN(
        n2507) );
  aoi22d1 U2749 ( .A1(n2337), .A2(n3233), .B1(pll_trim[0]), .B2(n2336), .ZN(
        n2506) );
  inv0d0 U2750 ( .I(n2339), .ZN(n2338) );
  aoi22d1 U2751 ( .A1(n2339), .A2(n3260), .B1(\gpio_configure[12][10] ), .B2(
        n2338), .ZN(n2505) );
  inv0d0 U2752 ( .I(n2535), .ZN(n2343) );
  aoi22d1 U2753 ( .A1(n2535), .A2(n3242), .B1(\gpio_configure[11][1] ), .B2(
        n2343), .ZN(n2504) );
  aoi22d1 U2754 ( .A1(n2535), .A2(n3233), .B1(\gpio_configure[11][0] ), .B2(
        n2343), .ZN(n2503) );
  aoi22d1 U2755 ( .A1(n3105), .A2(n3230), .B1(\gpio_configure[36][12] ), .B2(
        n3104), .ZN(n2502) );
  aoi22d1 U2756 ( .A1(n3105), .A2(n3231), .B1(\gpio_configure[36][11] ), .B2(
        n3104), .ZN(n2501) );
  aoi22d1 U2757 ( .A1(n3107), .A2(n3242), .B1(\gpio_configure[35][1] ), .B2(
        n3106), .ZN(n2500) );
  aoi22d1 U2758 ( .A1(n3107), .A2(n3233), .B1(\gpio_configure[35][0] ), .B2(
        n3106), .ZN(n2499) );
  aoi22d1 U2759 ( .A1(n3109), .A2(n3157), .B1(\gpio_configure[20][10] ), .B2(
        n3108), .ZN(n2498) );
  aoi22d1 U2760 ( .A1(n3111), .A2(n3242), .B1(\gpio_configure[19][1] ), .B2(
        n3110), .ZN(n2497) );
  aoi22d1 U2761 ( .A1(n3111), .A2(n3272), .B1(\gpio_configure[19][0] ), .B2(
        n3110), .ZN(n2496) );
  aoi22d1 U2762 ( .A1(n3113), .A2(n3204), .B1(\gpio_configure[24][10] ), .B2(
        n3112), .ZN(n2495) );
  aoi22d1 U2763 ( .A1(n3115), .A2(n3242), .B1(\gpio_configure[23][1] ), .B2(
        n3114), .ZN(n2494) );
  aoi22d1 U2764 ( .A1(n3115), .A2(n3272), .B1(\gpio_configure[23][0] ), .B2(
        n3114), .ZN(n2493) );
  aoi22d1 U2765 ( .A1(n3117), .A2(n3204), .B1(\gpio_configure[32][10] ), .B2(
        n3116), .ZN(n2492) );
  aoi22d1 U2766 ( .A1(n3119), .A2(n3242), .B1(\gpio_configure[31][1] ), .B2(
        n3118), .ZN(n2491) );
  aoi22d1 U2767 ( .A1(n3119), .A2(n3272), .B1(\gpio_configure[31][0] ), .B2(
        n3118), .ZN(n2490) );
  aoi22d1 U2768 ( .A1(n3121), .A2(n3260), .B1(\gpio_configure[28][10] ), .B2(
        n3120), .ZN(n2489) );
  aoi22d1 U2769 ( .A1(n3123), .A2(n3242), .B1(\gpio_configure[27][1] ), .B2(
        n3122), .ZN(n2488) );
  aoi22d1 U2770 ( .A1(n3123), .A2(n3272), .B1(\gpio_configure[27][0] ), .B2(
        n3122), .ZN(n2487) );
  inv0d0 U2771 ( .I(n3125), .ZN(n3124) );
  aoi22d1 U2772 ( .A1(n3125), .A2(n3204), .B1(\gpio_configure[11][10] ), .B2(
        n3124), .ZN(n2486) );
  aoi22d1 U2773 ( .A1(n3127), .A2(n3270), .B1(\gpio_configure[10][1] ), .B2(
        n3126), .ZN(n2485) );
  aoi22d1 U2774 ( .A1(n3127), .A2(n3272), .B1(\gpio_configure[10][0] ), .B2(
        n3126), .ZN(n2484) );
  inv0d0 U2775 ( .I(n3129), .ZN(n3128) );
  aoi22d1 U2776 ( .A1(n3129), .A2(n3204), .B1(pll_div[2]), .B2(n3128), .ZN(
        n2483) );
  inv0d0 U2777 ( .I(n3131), .ZN(n3130) );
  aoi22d1 U2778 ( .A1(n3131), .A2(n3231), .B1(\gpio_configure[3][11] ), .B2(
        n3130), .ZN(n2482) );
  inv0d0 U2779 ( .I(n3133), .ZN(n3132) );
  aoi22d1 U2780 ( .A1(n3133), .A2(n3204), .B1(\gpio_configure[7][10] ), .B2(
        n3132), .ZN(n2481) );
  inv0d0 U2781 ( .I(n3135), .ZN(n3134) );
  aoi22d1 U2782 ( .A1(n3135), .A2(n3270), .B1(\gpio_configure[6][1] ), .B2(
        n3134), .ZN(n2480) );
  aoi22d1 U2783 ( .A1(n3135), .A2(n3272), .B1(\gpio_configure[6][0] ), .B2(
        n3134), .ZN(n2479) );
  inv0d0 U2784 ( .I(n3137), .ZN(n3136) );
  aoi22d1 U2785 ( .A1(n3137), .A2(n3157), .B1(\gpio_configure[15][10] ), .B2(
        n3136), .ZN(n2478) );
  inv0d0 U2786 ( .I(n3139), .ZN(n3138) );
  aoi22d1 U2787 ( .A1(n3139), .A2(n3270), .B1(\gpio_configure[14][1] ), .B2(
        n3138), .ZN(n2477) );
  aoi22d1 U2788 ( .A1(n3139), .A2(n3233), .B1(\gpio_configure[14][0] ), .B2(
        n3138), .ZN(n2476) );
  aoi22d1 U2789 ( .A1(n3141), .A2(n3157), .B1(\gpio_configure[35][10] ), .B2(
        n3140), .ZN(n2475) );
  aoi22d1 U2790 ( .A1(n3143), .A2(n3270), .B1(\gpio_configure[34][1] ), .B2(
        n3142), .ZN(n2474) );
  aoi22d1 U2791 ( .A1(n3143), .A2(n3233), .B1(\gpio_configure[34][0] ), .B2(
        n3142), .ZN(n2473) );
  aoi22d1 U2792 ( .A1(n3145), .A2(n3157), .B1(\gpio_configure[19][10] ), .B2(
        n3144), .ZN(n2472) );
  inv0d0 U2793 ( .I(n3147), .ZN(n3146) );
  aoi22d1 U2794 ( .A1(n3147), .A2(n3270), .B1(\gpio_configure[18][1] ), .B2(
        n3146), .ZN(n2471) );
  aoi22d1 U2795 ( .A1(n3147), .A2(n3233), .B1(\gpio_configure[18][0] ), .B2(
        n3146), .ZN(n2470) );
  aoi22d1 U2796 ( .A1(n3149), .A2(n3157), .B1(\gpio_configure[23][10] ), .B2(
        n3148), .ZN(n2469) );
  inv0d0 U2797 ( .I(n3151), .ZN(n3150) );
  aoi22d1 U2798 ( .A1(n3151), .A2(n3270), .B1(\gpio_configure[22][1] ), .B2(
        n3150), .ZN(n2468) );
  aoi22d1 U2799 ( .A1(n3151), .A2(n3233), .B1(\gpio_configure[22][0] ), .B2(
        n3150), .ZN(n2467) );
  aoi22d1 U2800 ( .A1(n3153), .A2(n3157), .B1(\gpio_configure[31][10] ), .B2(
        n3152), .ZN(n2466) );
  aoi22d1 U2801 ( .A1(n3155), .A2(n3270), .B1(\gpio_configure[30][1] ), .B2(
        n3154), .ZN(n2465) );
  aoi22d1 U2802 ( .A1(n3155), .A2(n3268), .B1(\gpio_configure[30][0] ), .B2(
        n3154), .ZN(n2464) );
  aoi22d1 U2803 ( .A1(n3158), .A2(n3157), .B1(\gpio_configure[27][10] ), .B2(
        n3156), .ZN(n2463) );
  aoi22d1 U2804 ( .A1(n3160), .A2(n3270), .B1(\gpio_configure[26][1] ), .B2(
        n3159), .ZN(n2462) );
  aoi22d1 U2805 ( .A1(n3160), .A2(n3233), .B1(\gpio_configure[26][0] ), .B2(
        n3159), .ZN(n2461) );
  aoi22d1 U2806 ( .A1(n3162), .A2(n3260), .B1(\gpio_configure[14][10] ), .B2(
        n3161), .ZN(n2460) );
  inv0d0 U2807 ( .I(n3164), .ZN(n3163) );
  aoi22d1 U2808 ( .A1(n3164), .A2(n3242), .B1(\gpio_configure[13][1] ), .B2(
        n3163), .ZN(n2459) );
  aoi22d1 U2809 ( .A1(n3164), .A2(n3272), .B1(\gpio_configure[13][0] ), .B2(
        n3163), .ZN(n2458) );
  inv0d0 U2810 ( .I(n3166), .ZN(n3165) );
  aoi22d1 U2811 ( .A1(n3166), .A2(n3260), .B1(\gpio_configure[10][10] ), .B2(
        n3165), .ZN(n2457) );
  inv0d0 U2812 ( .I(n3168), .ZN(n3167) );
  aoi22d1 U2813 ( .A1(n3168), .A2(n3266), .B1(\gpio_configure[9][1] ), .B2(
        n3167), .ZN(n2456) );
  aoi22d1 U2814 ( .A1(n3168), .A2(n3233), .B1(\gpio_configure[9][0] ), .B2(
        n3167), .ZN(n2455) );
  nr02d0 U2815 ( .A1(n3170), .A2(n3169), .ZN(n3172) );
  inv0d0 U2816 ( .I(n3172), .ZN(n3171) );
  aoi22d1 U2817 ( .A1(n3172), .A2(n3266), .B1(pll_trim[25]), .B2(n3171), .ZN(
        n2454) );
  aoi22d1 U2818 ( .A1(n3172), .A2(n3272), .B1(pll_trim[24]), .B2(n3171), .ZN(
        n2453) );
  aoi22d1 U2819 ( .A1(n3174), .A2(n3266), .B1(pll_sel[1]), .B2(n3173), .ZN(
        n2452) );
  aoi22d1 U2820 ( .A1(n3174), .A2(n3230), .B1(pll90_sel[1]), .B2(n3173), .ZN(
        n2451) );
  inv0d0 U2821 ( .I(n3176), .ZN(n3175) );
  aoi22d1 U2822 ( .A1(n3176), .A2(n3204), .B1(\gpio_configure[6][10] ), .B2(
        n3175), .ZN(n2450) );
  inv0d0 U2823 ( .I(n3178), .ZN(n3177) );
  aoi22d1 U2824 ( .A1(n3178), .A2(n3266), .B1(\gpio_configure[5][1] ), .B2(
        n3177), .ZN(n2449) );
  aoi22d1 U2825 ( .A1(n3178), .A2(n3272), .B1(\gpio_configure[5][0] ), .B2(
        n3177), .ZN(n2448) );
  inv0d0 U2826 ( .I(n3180), .ZN(n3179) );
  aoi22d1 U2827 ( .A1(n3180), .A2(n3266), .B1(pll_dco_ena), .B2(n3179), .ZN(
        n2447) );
  nd02d0 U2828 ( .A1(n858), .A2(n3228), .ZN(n3182) );
  aoim22d1 U2829 ( .A1(pll_bypass), .A2(n3182), .B1(n3182), .B2(n3181), .Z(
        n2446) );
  inv0d0 U2830 ( .I(n3184), .ZN(n3183) );
  aoi22d1 U2831 ( .A1(n3184), .A2(n3204), .B1(\gpio_configure[2][10] ), .B2(
        n3183), .ZN(n2445) );
  aoi22d1 U2832 ( .A1(n3186), .A2(n3266), .B1(\gpio_configure[37][1] ), .B2(
        n3185), .ZN(n2444) );
  aoi22d1 U2833 ( .A1(n3186), .A2(n3272), .B1(\gpio_configure[37][0] ), .B2(
        n3185), .ZN(n2443) );
  aoi22d1 U2834 ( .A1(n3188), .A2(n3204), .B1(\gpio_configure[22][10] ), .B2(
        n3187), .ZN(n2442) );
  inv0d0 U2835 ( .I(n3190), .ZN(n3189) );
  aoi22d1 U2836 ( .A1(n3190), .A2(n3266), .B1(\gpio_configure[21][1] ), .B2(
        n3189), .ZN(n2441) );
  aoi22d1 U2837 ( .A1(n3190), .A2(n3272), .B1(\gpio_configure[21][0] ), .B2(
        n3189), .ZN(n2440) );
  aoi22d1 U2838 ( .A1(n3192), .A2(n3204), .B1(\gpio_configure[34][10] ), .B2(
        n3191), .ZN(n2439) );
  aoi22d1 U2839 ( .A1(n3194), .A2(n3270), .B1(\gpio_configure[33][1] ), .B2(
        n3193), .ZN(n2438) );
  aoi22d1 U2840 ( .A1(n3194), .A2(n3268), .B1(\gpio_configure[33][0] ), .B2(
        n3193), .ZN(n2437) );
  aoi22d1 U2841 ( .A1(n3196), .A2(n3204), .B1(\gpio_configure[18][10] ), .B2(
        n3195), .ZN(n2436) );
  inv0d0 U2842 ( .I(n3198), .ZN(n3197) );
  aoi22d1 U2843 ( .A1(n3198), .A2(n3270), .B1(\gpio_configure[17][1] ), .B2(
        n3197), .ZN(n2435) );
  aoi22d1 U2844 ( .A1(n3198), .A2(n3268), .B1(\gpio_configure[17][0] ), .B2(
        n3197), .ZN(n2434) );
  aoi22d1 U2845 ( .A1(n3200), .A2(n3204), .B1(\gpio_configure[30][10] ), .B2(
        n3199), .ZN(n2433) );
  aoi22d1 U2846 ( .A1(n3202), .A2(n3242), .B1(\gpio_configure[29][1] ), .B2(
        n3201), .ZN(n2432) );
  aoi22d1 U2847 ( .A1(n3202), .A2(n3268), .B1(\gpio_configure[29][0] ), .B2(
        n3201), .ZN(n2431) );
  aoi22d1 U2848 ( .A1(n3205), .A2(n3204), .B1(\gpio_configure[26][10] ), .B2(
        n3203), .ZN(n2430) );
  aoi22d1 U2849 ( .A1(n3207), .A2(n3266), .B1(\gpio_configure[25][1] ), .B2(
        n3206), .ZN(n2429) );
  aoi22d1 U2850 ( .A1(n3207), .A2(n3268), .B1(\gpio_configure[25][0] ), .B2(
        n3206), .ZN(n2428) );
  aoi22d1 U2851 ( .A1(n3209), .A2(n3260), .B1(\gpio_configure[5][10] ), .B2(
        n3208), .ZN(n2427) );
  inv0d0 U2852 ( .I(n3211), .ZN(n3210) );
  aoi22d1 U2853 ( .A1(n3211), .A2(n3270), .B1(\gpio_configure[4][1] ), .B2(
        n3210), .ZN(n2426) );
  aoi22d1 U2854 ( .A1(n3211), .A2(n3268), .B1(\gpio_configure[4][0] ), .B2(
        n3210), .ZN(n2425) );
  inv0d0 U2855 ( .I(n3213), .ZN(n3212) );
  aoi22d1 U2856 ( .A1(n3213), .A2(n3260), .B1(\gpio_configure[13][10] ), .B2(
        n3212), .ZN(n2424) );
  inv0d0 U2857 ( .I(n3215), .ZN(n3214) );
  aoi22d1 U2858 ( .A1(n3215), .A2(n3266), .B1(\gpio_configure[12][1] ), .B2(
        n3214), .ZN(n2423) );
  aoi22d1 U2859 ( .A1(n3215), .A2(n3272), .B1(\gpio_configure[12][0] ), .B2(
        n3214), .ZN(n2422) );
  inv0d0 U2860 ( .I(n3217), .ZN(n3216) );
  aoi22d1 U2861 ( .A1(n3217), .A2(n3260), .B1(\gpio_configure[17][10] ), .B2(
        n3216), .ZN(n2421) );
  inv0d0 U2862 ( .I(n3219), .ZN(n3218) );
  aoi22d1 U2863 ( .A1(n3219), .A2(n3242), .B1(\gpio_configure[16][1] ), .B2(
        n3218), .ZN(n2420) );
  aoi22d1 U2864 ( .A1(n3219), .A2(n3233), .B1(\gpio_configure[16][0] ), .B2(
        n3218), .ZN(n2419) );
  aoi22d1 U2865 ( .A1(n3221), .A2(n3230), .B1(\gpio_configure[1][12] ), .B2(
        n3220), .ZN(n2418) );
  aoi22d1 U2866 ( .A1(n3221), .A2(n3231), .B1(\gpio_configure[1][11] ), .B2(
        n3220), .ZN(n2417) );
  aoi22d1 U2867 ( .A1(n3223), .A2(n3270), .B1(\gpio_configure[0][1] ), .B2(
        n3222), .ZN(n2416) );
  aoi22d1 U2868 ( .A1(n3223), .A2(n3233), .B1(\gpio_configure[0][0] ), .B2(
        n3222), .ZN(n2415) );
  inv0d0 U2869 ( .I(n3225), .ZN(n3224) );
  aoi22d1 U2870 ( .A1(n3225), .A2(n3260), .B1(\gpio_configure[9][10] ), .B2(
        n3224), .ZN(n2414) );
  inv0d0 U2871 ( .I(n3227), .ZN(n3226) );
  aoi22d1 U2872 ( .A1(n3227), .A2(n3266), .B1(\gpio_configure[8][1] ), .B2(
        n3226), .ZN(n2413) );
  aoi22d1 U2873 ( .A1(n3227), .A2(n3272), .B1(\gpio_configure[8][0] ), .B2(
        n3226), .ZN(n2412) );
  nd02d0 U2874 ( .A1(n3229), .A2(n3228), .ZN(n3232) );
  inv0d0 U2875 ( .I(n3232), .ZN(n3234) );
  aoi22d1 U2876 ( .A1(n3234), .A2(n3235), .B1(pll_trim[23]), .B2(n3232), .ZN(
        n2411) );
  aoi22d1 U2877 ( .A1(n3234), .A2(n3236), .B1(pll_trim[22]), .B2(n3232), .ZN(
        n2410) );
  aoi22d1 U2878 ( .A1(n3234), .A2(n3237), .B1(pll_trim[21]), .B2(n3232), .ZN(
        n2409) );
  aoi22d1 U2879 ( .A1(n3234), .A2(n3230), .B1(pll_trim[20]), .B2(n3232), .ZN(
        n2408) );
  aoi22d1 U2880 ( .A1(n3234), .A2(n3231), .B1(pll_trim[19]), .B2(n3232), .ZN(
        n2407) );
  aoi22d1 U2881 ( .A1(n3234), .A2(n3260), .B1(pll_trim[18]), .B2(n3232), .ZN(
        n2406) );
  aoi22d1 U2882 ( .A1(n3234), .A2(n3266), .B1(pll_trim[17]), .B2(n3232), .ZN(
        n2405) );
  aoi22d1 U2883 ( .A1(n3234), .A2(n3233), .B1(pll_trim[16]), .B2(n3232), .ZN(
        n2404) );
  inv0d0 U2884 ( .I(n3239), .ZN(n3238) );
  aoi22d1 U2885 ( .A1(n3239), .A2(n3235), .B1(pll_trim[15]), .B2(n3238), .ZN(
        n2403) );
  aoi22d1 U2886 ( .A1(n3239), .A2(n3236), .B1(pll_trim[14]), .B2(n3238), .ZN(
        n2402) );
  aoi22d1 U2887 ( .A1(n3239), .A2(n3237), .B1(pll_trim[13]), .B2(n3238), .ZN(
        n2401) );
  aoi22d1 U2888 ( .A1(n3239), .A2(n3247), .B1(pll_trim[11]), .B2(n3238), .ZN(
        n2400) );
  aoi22d1 U2889 ( .A1(n3239), .A2(n3260), .B1(pll_trim[10]), .B2(n3238), .ZN(
        n2399) );
  aoi22d1 U2890 ( .A1(n3239), .A2(n3266), .B1(pll_trim[9]), .B2(n3238), .ZN(
        n2398) );
  aoi22d1 U2891 ( .A1(n3239), .A2(n3268), .B1(pll_trim[8]), .B2(n3238), .ZN(
        n2397) );
  aoi22d1 U2892 ( .A1(n3241), .A2(n3260), .B1(\gpio_configure[25][10] ), .B2(
        n3240), .ZN(n2396) );
  aoi22d1 U2893 ( .A1(n3244), .A2(n3242), .B1(\gpio_configure[24][1] ), .B2(
        n3243), .ZN(n2395) );
  aoi22d1 U2894 ( .A1(n3244), .A2(n3268), .B1(\gpio_configure[24][0] ), .B2(
        n3243), .ZN(n2394) );
  aoi22d1 U2895 ( .A1(n3248), .A2(n3245), .B1(\gpio_configure[37][12] ), .B2(
        n3246), .ZN(n2393) );
  aoi22d1 U2896 ( .A1(n3248), .A2(n3247), .B1(\gpio_configure[37][11] ), .B2(
        n3246), .ZN(n2392) );
  aoi22d1 U2897 ( .A1(n3250), .A2(n3266), .B1(\gpio_configure[36][1] ), .B2(
        n3249), .ZN(n2391) );
  aoi22d1 U2898 ( .A1(n3250), .A2(n3268), .B1(\gpio_configure[36][0] ), .B2(
        n3249), .ZN(n2390) );
  aoi22d1 U2899 ( .A1(n3252), .A2(n3260), .B1(\gpio_configure[21][10] ), .B2(
        n3251), .ZN(n2389) );
  inv0d0 U2900 ( .I(n3254), .ZN(n3253) );
  aoi22d1 U2901 ( .A1(n3254), .A2(n3270), .B1(\gpio_configure[20][1] ), .B2(
        n3253), .ZN(n2388) );
  aoi22d1 U2902 ( .A1(n3254), .A2(n3268), .B1(\gpio_configure[20][0] ), .B2(
        n3253), .ZN(n2387) );
  aoi22d1 U2903 ( .A1(n3256), .A2(n3260), .B1(\gpio_configure[33][10] ), .B2(
        n3255), .ZN(n2386) );
  aoi22d1 U2904 ( .A1(n3258), .A2(n3266), .B1(\gpio_configure[32][1] ), .B2(
        n3257), .ZN(n2385) );
  aoi22d1 U2905 ( .A1(n3258), .A2(n3268), .B1(\gpio_configure[32][0] ), .B2(
        n3257), .ZN(n2384) );
  aoi22d1 U2906 ( .A1(n3261), .A2(n3260), .B1(\gpio_configure[29][10] ), .B2(
        n3259), .ZN(n2383) );
  aoi22d1 U2907 ( .A1(n3263), .A2(n3270), .B1(\gpio_configure[28][1] ), .B2(
        n3262), .ZN(n2382) );
  aoi22d1 U2908 ( .A1(n3263), .A2(n3268), .B1(\gpio_configure[28][0] ), .B2(
        n3262), .ZN(n2381) );
  inv0d0 U2909 ( .I(n3265), .ZN(n3264) );
  aoi22d1 U2910 ( .A1(n3265), .A2(n3268), .B1(\gpio_configure[3][0] ), .B2(
        n3264), .ZN(n2380) );
  aoi22d1 U2911 ( .A1(n3269), .A2(n3266), .B1(\gpio_configure[2][1] ), .B2(
        n3267), .ZN(n2379) );
  aoi22d1 U2912 ( .A1(n3269), .A2(n3268), .B1(\gpio_configure[2][0] ), .B2(
        n3267), .ZN(n2378) );
  aoi22d1 U2913 ( .A1(n3273), .A2(n3270), .B1(\gpio_configure[1][1] ), .B2(
        n3271), .ZN(n2377) );
  aoi22d1 U2914 ( .A1(n3273), .A2(n3272), .B1(\gpio_configure[1][0] ), .B2(
        n3271), .ZN(n2376) );
  nd03d0 U2915 ( .A1(wbbd_state[1]), .A2(n3274), .A3(n3292), .ZN(n3276) );
  nr02d1 U2916 ( .A1(wbbd_state[2]), .A2(n3276), .ZN(n3286) );
  aoim22d1 U2917 ( .A1(n3286), .A2(n3279), .B1(wb_dat_o[7]), .B2(n3286), .Z(
        n2375) );
  nr04d2 U2918 ( .A1(wb_rstn_i), .A2(wbbd_state[1]), .A3(n3277), .A4(n3275), 
        .ZN(n3287) );
  aoim22d1 U2919 ( .A1(n3287), .A2(n3279), .B1(wb_dat_o[15]), .B2(n3287), .Z(
        n2374) );
  nr02d1 U2920 ( .A1(n3277), .A2(n3276), .ZN(n3288) );
  aoim22d1 U2921 ( .A1(n3288), .A2(n3279), .B1(wb_dat_o[23]), .B2(n3288), .Z(
        n2373) );
  nr02d1 U2922 ( .A1(wb_rstn_i), .A2(n3278), .ZN(n3290) );
  aoim22d1 U2923 ( .A1(n3290), .A2(n3279), .B1(wb_dat_o[31]), .B2(n3290), .Z(
        n2372) );
  aoim22d1 U2924 ( .A1(n3286), .A2(n3280), .B1(wb_dat_o[4]), .B2(n3286), .Z(
        n2371) );
  aoim22d1 U2925 ( .A1(n3287), .A2(n3280), .B1(wb_dat_o[12]), .B2(n3287), .Z(
        n2370) );
  aoim22d1 U2926 ( .A1(n3288), .A2(n3280), .B1(wb_dat_o[20]), .B2(n3288), .Z(
        n2369) );
  aoim22d1 U2927 ( .A1(n3290), .A2(n3280), .B1(wb_dat_o[28]), .B2(n3290), .Z(
        n2368) );
  aoim22d1 U2928 ( .A1(n3286), .A2(n3281), .B1(wb_dat_o[5]), .B2(n3286), .Z(
        n2367) );
  aoim22d1 U2929 ( .A1(n3287), .A2(n3281), .B1(wb_dat_o[13]), .B2(n3287), .Z(
        n2366) );
  aoim22d1 U2930 ( .A1(n3288), .A2(n3281), .B1(wb_dat_o[21]), .B2(n3288), .Z(
        n2365) );
  aoim22d1 U2931 ( .A1(n3290), .A2(n3281), .B1(wb_dat_o[29]), .B2(n3290), .Z(
        n2364) );
  aoim22d1 U2932 ( .A1(n3286), .A2(n3282), .B1(wb_dat_o[6]), .B2(n3286), .Z(
        n2363) );
  aoim22d1 U2933 ( .A1(n3287), .A2(n3282), .B1(wb_dat_o[14]), .B2(n3287), .Z(
        n2362) );
  aoim22d1 U2934 ( .A1(n3288), .A2(n3282), .B1(wb_dat_o[22]), .B2(n3288), .Z(
        n2361) );
  aoim22d1 U2935 ( .A1(n3290), .A2(n3282), .B1(wb_dat_o[30]), .B2(n3290), .Z(
        n2360) );
  aoim22d1 U2936 ( .A1(n3286), .A2(n3283), .B1(wb_dat_o[0]), .B2(n3286), .Z(
        n2359) );
  aoim22d1 U2937 ( .A1(n3287), .A2(n3283), .B1(wb_dat_o[8]), .B2(n3287), .Z(
        n2358) );
  aoim22d1 U2938 ( .A1(n3288), .A2(n3283), .B1(wb_dat_o[16]), .B2(n3288), .Z(
        n2357) );
  aoim22d1 U2939 ( .A1(n3290), .A2(n3283), .B1(wb_dat_o[24]), .B2(n3290), .Z(
        n2356) );
  aoim22d1 U2940 ( .A1(n3286), .A2(n3284), .B1(wb_dat_o[3]), .B2(n3286), .Z(
        n2355) );
  aoim22d1 U2941 ( .A1(n3287), .A2(n3284), .B1(wb_dat_o[11]), .B2(n3287), .Z(
        n2354) );
  aoim22d1 U2942 ( .A1(n3288), .A2(n3284), .B1(wb_dat_o[19]), .B2(n3288), .Z(
        n2353) );
  aoim22d1 U2943 ( .A1(n3290), .A2(n3284), .B1(wb_dat_o[27]), .B2(n3290), .Z(
        n2352) );
  aoim22d1 U2944 ( .A1(n3286), .A2(n3285), .B1(wb_dat_o[2]), .B2(n3286), .Z(
        n2351) );
  aoim22d1 U2945 ( .A1(n3287), .A2(n3285), .B1(wb_dat_o[10]), .B2(n3287), .Z(
        n2350) );
  aoim22d1 U2946 ( .A1(n3288), .A2(n3285), .B1(wb_dat_o[18]), .B2(n3288), .Z(
        n2349) );
  aoim22d1 U2947 ( .A1(n3290), .A2(n3285), .B1(wb_dat_o[26]), .B2(n3290), .Z(
        n2348) );
  aoim22d1 U2948 ( .A1(n3286), .A2(n3289), .B1(wb_dat_o[1]), .B2(n3286), .Z(
        n2347) );
  aoim22d1 U2949 ( .A1(n3287), .A2(n3289), .B1(wb_dat_o[9]), .B2(n3287), .Z(
        n2346) );
  aoim22d1 U2950 ( .A1(n3288), .A2(n3289), .B1(wb_dat_o[17]), .B2(n3288), .Z(
        n2345) );
  aoim22d1 U2951 ( .A1(n3290), .A2(n3289), .B1(wb_dat_o[25]), .B2(n3290), .Z(
        n2344) );
endmodule


